module top( V32(0), V32(1), V32(2), V32(3), V56(0), V289(0), V10(0), V13(0), V35(0), V203(0), V288(6), V288(7), V248(0), V249(0), V62(0), V59(0), V174(0), V215(0), V66(0), V70(0), V43(0), V214(0), V37(0), V271(0), V40(0), V45(0), V149(7), V149(6), V149(5), V149(4), V1(0), V7(0), V34(0), V243(0), V244(0), V245(0), V246(0), V247(0), V293(0), V302(0), V270(0), V269(0), V274(0), V202(0), V275(0), V257(7), V257(5), V257(3), V257(1), V257(2), V257(4), V257(6), V9(0), V149(0), V149(1), V149(2), V149(3), V169(1), V165(0), V165(2), V165(4), V165(5), V165(6), V165(7), V165(1), V88(2), V88(3), V55(0), V169(0), V52(0), V5(0), V6(0), V12(0), V11(0), V4(0), V165(3), V51(0), V65(0), V290(0), V279(0), V280(0), V288(4), V288(2), V288(0), V258(0), V229(5), V229(4), V229(3), V229(2), V229(1), V229(0), V223(5), V223(4), V223(3), V223(2), V223(1), V223(0), V189(5), V189(4), V189(3), V189(2), V189(1), V189(0), V183(5), V183(4), V183(3), V183(2), V183(1), V183(0), V239(4), V239(3), V239(2), V239(1), V239(0), V234(4), V234(3), V234(2), V234(1), V234(0), V199(4), V199(3), V199(2), V199(1), V199(0), V194(4), V194(3), V194(2), V194(1), V194(0), V257(0), V32(8), V32(7), V32(6), V32(5), V32(4), V32(11), V32(10), V32(9), V88(1), V88(0), V84(5), V84(4), V84(3), V84(2), V84(1), V84(0), V78(5), V78(4), V2(0), V3(0), V14(0), V213(0), V213(5), V213(4), V213(3), V213(2), V213(1), V268(5), V268(3), V268(1), V268(2), V268(4), V8(0), V60(0), V53(0), V57(0), V109(0), V277(0), V278(0), V259(0), V260(0), V67(0), V68(0), V69(0), V216(0), V175(0), V177(0), V172(0), V171(0), V50(0), V63(0), V71(0), V292(0), V291(0), V91(0), V91(1), V294(0), V207(0), V295(0), V204(0), V205(0), V261(0), V262(0), V100(0), V100(5), V100(4), V100(3), V100(2), V100(1), V240(0), V242(0), V241(0), V33(0), V16(0), V15(0), V101(0), V268(0), V288(1), V288(3), V288(5), V301(0), V108(0), V108(1), V108(2), V108(3), V108(4), V108(5), V124(5), V124(4), V124(3), V124(2), V124(1), V124(0), V132(7), V132(6), V132(5), V132(4), V132(3), V132(2), V132(1), V132(0), V118(5), V118(4), V118(3), V118(2), V118(1), V118(0), V118(7), V118(6), V46(0), V48(0), V102(0), V110(0), V134(1), V134(0), V272(0), V78(2), V78(3), V39(0), V38(0), V42(0), V44(0), V41(0), V78(1), V78(0), V94(0), V94(1), V321(2), V356, V357, V373, V375(0), V377, V393(0), V398(0), V410(0), V423(0), V432, V435(0), V500(0), V508(0), V511(0), V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, V572(9), V572(8), V572(7), V572(6), V572(5), V572(4), V572(3), V572(2), V572(1), V572(0), V585(0), V587, V591(0), V597(0), V603(0), V609(0), V620, V621, V630, V634(0), V640(0), V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V798(0), V801, V802(0), V821(0), V826(0), V966, V986, V1213(11), V1213(10), V1213(9), V1213(8), V1213(7), V1213(6), V1213(5), V1213(4), V1213(3), V1213(2), V1213(1), V1213(0), V1243(9), V1243(8), V1243(7), V1243(6), V1243(5), V1243(4), V1243(3), V1243(2), V1243(1), V1243(0), V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, V1274(0), V1281(0), V1297(4), V1297(3), V1297(2), V1297(1), V1297(0), V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1392(0), V1423, V1426, V1428, V1429, V1431, V1432, V1439(0), V1440(0), V1451(0), V1459(0), V1467(0), V1470, V1480(0), V1481(0), V1492(0), V1495(0), V1512(3), V1512(2), V1512(1), V1536(0), V1537, V1539, V1552(1), V1552(0), V1613(0), V1613(1), V1620(0), V1629(0), V1645(0), V1652(0), V1669, V1671(0), V1679(0), V1693(0), V1709(4), V1709(3), V1709(2), V1709(1), V1709(0), V1717(0), V1719, V1726(0), V1736, V1741(0), V1745(0), V1757(0), V1758(0), V1759(0), V1760(0), V1771(1), V1771(0), V1781(1), V1781(0), V1829(9), V1829(8), V1829(7), V1829(6), V1829(5), V1829(4), V1829(3), V1829(2), V1829(1), V1829(0), V1832, V1833(0), V1863(0), V1864(0), V1896(0), V1897(0), V1898(0), V1899(0), V1900(0), V1901(0), V1921(5), V1921(4), V1921(3), V1921(2), V1921(1), V1921(0), V1953(1), V1953(7), V1953(6), V1953(5), V1953(4), V1953(3), V1953(2), V1953(0), V1960(1), V1960(0), V1968(0), V1992(1), V1992(0), V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374 );
  input V32(0), V32(1), V32(2), V32(3), V56(0), V289(0), V10(0), V13(0), V35(0), V203(0), V288(6), V288(7), V248(0), V249(0), V62(0), V59(0), V174(0), V215(0), V66(0), V70(0), V43(0), V214(0), V37(0), V271(0), V40(0), V45(0), V149(7), V149(6), V149(5), V149(4), V1(0), V7(0), V34(0), V243(0), V244(0), V245(0), V246(0), V247(0), V293(0), V302(0), V270(0), V269(0), V274(0), V202(0), V275(0), V257(7), V257(5), V257(3), V257(1), V257(2), V257(4), V257(6), V9(0), V149(0), V149(1), V149(2), V149(3), V169(1), V165(0), V165(2), V165(4), V165(5), V165(6), V165(7), V165(1), V88(2), V88(3), V55(0), V169(0), V52(0), V5(0), V6(0), V12(0), V11(0), V4(0), V165(3), V51(0), V65(0), V290(0), V279(0), V280(0), V288(4), V288(2), V288(0), V258(0), V229(5), V229(4), V229(3), V229(2), V229(1), V229(0), V223(5), V223(4), V223(3), V223(2), V223(1), V223(0), V189(5), V189(4), V189(3), V189(2), V189(1), V189(0), V183(5), V183(4), V183(3), V183(2), V183(1), V183(0), V239(4), V239(3), V239(2), V239(1), V239(0), V234(4), V234(3), V234(2), V234(1), V234(0), V199(4), V199(3), V199(2), V199(1), V199(0), V194(4), V194(3), V194(2), V194(1), V194(0), V257(0), V32(8), V32(7), V32(6), V32(5), V32(4), V32(11), V32(10), V32(9), V88(1), V88(0), V84(5), V84(4), V84(3), V84(2), V84(1), V84(0), V78(5), V78(4), V2(0), V3(0), V14(0), V213(0), V213(5), V213(4), V213(3), V213(2), V213(1), V268(5), V268(3), V268(1), V268(2), V268(4), V8(0), V60(0), V53(0), V57(0), V109(0), V277(0), V278(0), V259(0), V260(0), V67(0), V68(0), V69(0), V216(0), V175(0), V177(0), V172(0), V171(0), V50(0), V63(0), V71(0), V292(0), V291(0), V91(0), V91(1), V294(0), V207(0), V295(0), V204(0), V205(0), V261(0), V262(0), V100(0), V100(5), V100(4), V100(3), V100(2), V100(1), V240(0), V242(0), V241(0), V33(0), V16(0), V15(0), V101(0), V268(0), V288(1), V288(3), V288(5), V301(0), V108(0), V108(1), V108(2), V108(3), V108(4), V108(5), V124(5), V124(4), V124(3), V124(2), V124(1), V124(0), V132(7), V132(6), V132(5), V132(4), V132(3), V132(2), V132(1), V132(0), V118(5), V118(4), V118(3), V118(2), V118(1), V118(0), V118(7), V118(6), V46(0), V48(0), V102(0), V110(0), V134(1), V134(0), V272(0), V78(2), V78(3), V39(0), V38(0), V42(0), V44(0), V41(0), V78(1), V78(0), V94(0), V94(1);
  output V321(2), V356, V357, V373, V375(0), V377, V393(0), V398(0), V410(0), V423(0), V432, V435(0), V500(0), V508(0), V511(0), V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, V572(9), V572(8), V572(7), V572(6), V572(5), V572(4), V572(3), V572(2), V572(1), V572(0), V585(0), V587, V591(0), V597(0), V603(0), V609(0), V620, V621, V630, V634(0), V640(0), V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, V798(0), V801, V802(0), V821(0), V826(0), V966, V986, V1213(11), V1213(10), V1213(9), V1213(8), V1213(7), V1213(6), V1213(5), V1213(4), V1213(3), V1213(2), V1213(1), V1213(0), V1243(9), V1243(8), V1243(7), V1243(6), V1243(5), V1243(4), V1243(3), V1243(2), V1243(1), V1243(0), V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, V1274(0), V1281(0), V1297(4), V1297(3), V1297(2), V1297(1), V1297(0), V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, V1392(0), V1423, V1426, V1428, V1429, V1431, V1432, V1439(0), V1440(0), V1451(0), V1459(0), V1467(0), V1470, V1480(0), V1481(0), V1492(0), V1495(0), V1512(3), V1512(2), V1512(1), V1536(0), V1537, V1539, V1552(1), V1552(0), V1613(0), V1613(1), V1620(0), V1629(0), V1645(0), V1652(0), V1669, V1671(0), V1679(0), V1693(0), V1709(4), V1709(3), V1709(2), V1709(1), V1709(0), V1717(0), V1719, V1726(0), V1736, V1741(0), V1745(0), V1757(0), V1758(0), V1759(0), V1760(0), V1771(1), V1771(0), V1781(1), V1781(0), V1829(9), V1829(8), V1829(7), V1829(6), V1829(5), V1829(4), V1829(3), V1829(2), V1829(1), V1829(0), V1832, V1833(0), V1863(0), V1864(0), V1896(0), V1897(0), V1898(0), V1899(0), V1900(0), V1901(0), V1921(5), V1921(4), V1921(3), V1921(2), V1921(1), V1921(0), V1953(1), V1953(7), V1953(6), V1953(5), V1953(4), V1953(3), V1953(2), V1953(0), V1960(1), V1960(0), V1968(0), V1992(1), V1992(0), V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374;
wire n485, n487, n489, n492, n493, n494, n497, n499, n500, n501, n3159, n509, n513, n3163, n523, n3173, n533, n534, n537, n538, n540, n542, n544, n545, n549, n552, n557, n565, n566, n567, n3186, n577, n578, n583, n587, n591, n593, n596, n598, n599, n626, n627, n628, n630, n631, n647, n651, n3201, n3208, n661, n667, n671, n673, n675, n676, n681, n684, n687, n690, n703, n3222, n713, n717, n727, n734, n740, n741, n747, n760, n766, n772, n782, n795, n809, n814, n3232, n823, n834, n842, n850, n857, n863, n869, n874, n3242, n883, n898, n3252, n907, n912, n3259, n916, n946, n960, n970, n976, n982, n992, n3266, n1001, n1022, n1055, n3276, n3275, n3274, n1086, n3282, n3289, n3291, n1114, n3298, n1131, n3305, n1148, n3314, n3325, n1173, n3330, n1190, n3338, n3337, n3336, n1207, n1212, n3351, n3352, n1235, n3358, n1252, n3367, n1269, n3372, n3381, n3380, n1304, n1307, n1309, n1311, n1313, n1321, n1329, n1334, n3403, n3404, n1344, n3412, n1358, n1363, n3420, n1377, n1382, n3428, n1396, n1401, n1406, n1407, n1408, n3438, n1414, n1420, n1421, n1426, n1429, n1431, n1435, n3447, n1443, n3451, n3450, n1454, n1457, n3466, n3465, n3474, n1476, n3479, n3486, n1500, n1504, n1510, n1511, n1513, n1514, n1518, n3495, n1523, n1541, n1547, n1565, n1571, n1576, n1579, n1580, n1584, n1586, n3501, n3510, n3509, n1601, n1604, n1608, n3523, n1616, n1620, n1621, n1626, n1628, n3535, n3540, n3539, n1668, n1672, n1679, n1688, n1692, n1702, n1711, n1715, n1725, n1734, n1738, n1745, n1751, n1760, n1764, n1771, n1777, n1786, n1790, n1797, n1803, n1812, n1816, n1822, n1830, n1836, n1840, n1846, n1854, n1858, n1860, n1864, n1865, n3631, n3638, n1903, n1912, n1915, n1920, n3650, n1937, n1946, n1949, n1954, n3666, n1972, n1981, n1984, n1989, n1998, n2012, n2020, n3694, n2029, n2038, n2043, n3701, n2059, n2067, n3718, n2076, n2085, n2090, n3725, n3732, n3733, n2115, n3742, n2124, n2133, n2138, n3749, n3753, n3758, n3775, n2207, n2213, n2216, n2219, n2221, n3791, n2225, n2228, n3799, n2233, n3802, n3808, n3810, n2251, n2254, n2259, n2261, n2263, n2266, n2277, n2278, n2286, n2298, n2301, n2306, n2307, n2308, n3829, n2314, n2317, n2320, n2328, n2336, n3837, n3851, n2366, n2369, n2380, n3868, n2397, n2402, n3887, n3886, n2413, n3897, n2424, n3901, n2429, n2430, n2439, n3911, n3922, n3927, n2508, n2509, n3942, n2535, n3956, n3962, n3965, n2585, n2591, n3979, n2603, n3988, n3997, n2657, n4010, n2671, n4018, n4017, n2690, n4024, n4023, n4030, n4029, n2734, n4036, n4035, n4042, n4041, n2775, n2778, n2781, n2789, n2794, n2797, n2804, n2811, n2824, n2831, n2841, n2848, n2851, n2867, n4069, n2884, n4075, n2892, n2897, n4084, n2911, n2915, n2917, n4102, n2975, n4109, n3056, n4116, n3102, n3103 ; 
assign n485 = ((((n30)*(~(n54)))*(n55))*(n56))*(~(n57)) ;
assign n487 = ((~(n54))*(~(n55)))*(~(n56)) ;
assign n489 = ((~(n54))*(n55))*(~(n56)) ;
assign n492 = (((((~(n54))*(n55))*(~(n56)))*(n27))*(n29))*(~(n57)) ;
assign n493 = (n30)*((((n27)*(n29))*(~(n57)))*(n489)) ;
assign n494 = (n28)*((n30)*((((n27)*(n29))*(~(n57)))*(n489))) ;
assign n497 = (((((~(n54))*(n55))*(~(n56)))*(~(n27)))*(n29))*(~(n57)) ;
assign n499 = (((((~(n27))*(n29))*(~(n57)))*(n489))*(n28))*(n30) ;
assign n500 = (~((n28)*((n30)*((((n27)*(n29))*(~(n57)))*(n489)))))*(~((((((~(n27))*(n29))*(~(n57)))*(n489))*(n28))*(n30))) ;
assign n501 = (~(n70))*(~(n77)) ;
assign n3159 = (~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n68))*(~(n500)))*(n501))) ;
assign n509 = ((((n20)*(~(n61)))*(~(n62)))*(~(n63)))*(n76) ;
assign n513 = ((((~((~(n485))*(n3159)))*(n69))*(~(n183)))*(~(n184)))*(~(n509)) ;
assign n3163 = (((((n20)*(n62))*(n64))*(n192))*(n59))*(n60) ;
assign n523 = (((((n61)*(n63))*(n65))*(n76))*(n513))*(n3163) ;
assign n3173 = (((((n62)*(n63))*(n64))*(n59))*(n60))*(n61) ;
assign n533 = (~(n523))*(~(((((n65)*(n76))*(~(n190)))*(n192))*(n3173))) ;
assign n534 = (~(n193))*(n533) ;
assign n537 = (((~(n54))*(n55))*(n56))*(n57) ;
assign n538 = (~(n17))*(((((n30)*(~(n54)))*(n55))*(n56))*(~(n57))) ;
assign n540 = (n169)*(~((n168)*((~(n17))*(n485)))) ;
assign n542 = (~(n16))*(((((~(n54))*(n55))*(n56))*(n57))*(~(n540))) ;
assign n544 = ((~(n54))*(~(n55)))*(n56) ;
assign n545 = (~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56))) ;
assign n549 = ((((~(n30))*(~(n54)))*(n55))*(n56))*(~(n57)) ;
assign n552 = (~(n17))*(~(((~((~(n17))*(((((n30)*(~(n54)))*(n55))*(n56))*(~(n57)))))*(~(((((~(n30))*(~(n54)))*(n55))*(n56))*(~(n57)))))*((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56)))))) ;
assign n557 = ((~(((n537)*(~(n540)))*(~((~(n16))*(~(n164))))))*(~((n537)*(n540))))*(~(n552)) ;
assign n565 = (((((~(n16))*(n30))*(n534))*(n537))*(~(n540)))*(n557) ;
assign n566 = (~((((~(n54))*(n55))*(n56))*(n57)))*(~((~(n17))*(((((n30)*(~(n54)))*(n55))*(n56))*(~(n57))))) ;
assign n567 = (~(((((~(n30))*(~(n54)))*(n55))*(n56))*(~(n57))))*((~((((~(n54))*(n55))*(n56))*(n57)))*(~((~(n17))*(((((n30)*(~(n54)))*(n55))*(n56))*(~(n57)))))) ;
assign n3186 = (~((~(((~((~(n487))*(~(n544))))*(n119))*(n567)))*(~((((~(n487))*(~(n544)))*(n129))*(~(n567))))))*(n534) ;
assign n577 = ((~((((n46)*(~(n534)))*(~(n542)))*(n557)))*(~(((~(n542))*(~(n557)))*(n3186))))*(~(n565)) ;
assign n578 = (n513)*((~(n193))*(n533)) ;
assign n583 = (n513)*(~(((~(n5))*(~(n16)))*(~(n164)))) ;
assign n587 = (~((n3)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n134)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n591 = (n57)*(((~(n54))*(~(n55)))*(n56)) ;
assign n593 = (n164)*(~((~((~(n17))*(n485)))*(~((n57)*(n544))))) ;
assign n596 = ((((~(n54))*(n55))*(~(n56)))*((n27)*(~(n29))))*(~(n57)) ;
assign n598 = (n28)*((n30)*((((n27)*(~(n29)))*(~(n57)))*(n489))) ;
assign n599 = (~(n17))*(((~(n54))*(~(n55)))*(~(n56))) ;
assign n626 = (((((((~((~(n67))*((n66)*((((n29)*(~(n30)))*(~(n57)))*(n599)))))*(~((~(n67))*((~(n66))*((((n29)*(~(n30)))*(~(n57)))*(n599))))))*(~((~(n67))*((n66)*((((~(n57))*(n599))*(~(n29)))*(~(n30)))))))*(~((n67)*((~(n66))*((((~(n57))*(n599))*(~(n29)))*(~(n30)))))))*(~((n67)*((n66)*((((~(n57))*(n599))*(~(n29)))*(~(n30)))))))*(~((n67)*((~(n66))*((((n29)*(~(n30)))*(~(n57)))*(n599))))))*(~((((~(n57))*(n599))*(n29))*(n30))))*(~((((~(n57))*(n599))*(~(n29)))*(n30))) ;
assign n627 = (n58)*(~((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56))))) ;
assign n628 = (~(n626))*((n58)*(~((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56)))))) ;
assign n630 = (n57)*((~(n17))*(((~(n54))*(~(n55)))*(~(n56)))) ;
assign n631 = ((n58)*(~((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56))))))*((n57)*((~(n17))*(((~(n54))*(~(n55)))*(~(n56))))) ;
assign n647 = ((~((n30)*(((((~(n54))*(~(n55)))*(n56))*(~(n29)))*(~(n57)))))*(~((~(n30))*(((((~(n54))*(~(n55)))*(n56))*(~(n29)))*(~(n57))))))*(~((~(n30))*(((((~(n54))*(~(n55)))*(n56))*(n29))*(~(n57))))) ;
assign n651 = (((~((n538)*(~(n540))))*((~(n591))*(n626)))*(~(n630)))*(n647) ;
assign n3201 = (((~((n164)*((n627)*((n57)*(n599)))))*(~((n5)*((n627)*((n57)*(n599))))))*(~((n164)*((~(n626))*(n627)))))*(~((n5)*((~(n626))*(n627)))) ;
assign n3208 = (~(((~(((~(n5))*(~(n165)))*(~(n166))))*(~(n651)))*(n3201)))*(~(n598)) ;
assign n661 = (~(((((~(n5))*(n165))*(n534))*(~(n537)))*(~(n549))))*(n3208) ;
assign n667 = (~(((~((~((~(n578))*((~(n577))*(~(n578)))))*(~((n578)*((n578)*(~(n587)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n148))*(~(n661)))) ;
assign n671 = ((((~(n27))*(~(n29)))*(~(n30)))*(n57))*(n489) ;
assign n673 = ((~(n70))*(~(n77)))*((~(n28))*(n671)) ;
assign n675 = (~(n84))*(n208) ;
assign n676 = (~(n83))*(n209) ;
assign n681 = (~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))) ;
assign n684 = (~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))) ;
assign n687 = (~(((~(n84))*(n208))*((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681)))))))) ;
assign n690 = (n84)*(~(n208)) ;
assign n703 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n94)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n106))) ;
assign n3222 = (((~((~(n16))*((n537)*(~(n540)))))*((~(n557))*(~((n513)*(n534)))))*(~((n513)*(n534))))*(n534) ;
assign n713 = (~((((~((~(n593))*(~(n661))))*(n661))*(~(n703)))*(n3222)))*(~((((~(n593))*(~(n661)))*(n4))*(~(n661)))) ;
assign n717 = (n83)*(~(n209)) ;
assign n727 = (~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))) ;
assign n734 = (~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))) ;
assign n740 = ((~(((n84)*(~(n208)))*(~((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681)))))))))*(~((~((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681)))))))*(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))))) ;
assign n741 = (n84)*(n208) ;
assign n747 = (n83)*(n209) ;
assign n760 = (~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))) ;
assign n766 = (~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))) ;
assign n772 = (~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))) ;
assign n782 = (~((~(((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681)))))))))))))*(~((((~(n84))*(n208))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681)))))))*((~(((n84)*(~(n208)))*((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681))))))))*(~((~((n84)*(~(n208))))*(~((~((~((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727))))))*(~(((~(n83))*(n209))*(~(n681))))))*(~(((~(((n83)*(~(n209)))*(n727)))*(~((~((n83)*(~(n209))))*(~(n727)))))*(((~(n83))*(n209))*(~(n681)))))))))))) ;
assign n795 = (~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))*(~(((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))) ;
assign n809 = (~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~((~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))*(~(((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))))))))*(~(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))))))))*(~(((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))*(~(((~((~((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~(((~((~(((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734))))))*((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))*(~((((~((~(n734))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~(((n84)*(~(n208)))*(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~(((n84)*(~(n208)))*(~(n734)))))*(~((~(((n84)*(n208))*(n766)))*(~((~((n84)*(n208)))*(~(n766)))))))))*(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))))*(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))))))))))))))) ;
assign n814 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n96)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n108))) ;
assign n3232 = (((~((~(n16))*((n537)*(~(n540)))))*((~(n557))*(~((n513)*(n534)))))*(~((n513)*(n534))))*(n534) ;
assign n823 = (~((((~((~(n593))*(~(n661))))*(n661))*(~(n814)))*(n3232)))*(~((((~(n593))*(~(n661)))*(n2))*(~(n661)))) ;
assign n834 = (~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))) ;
assign n842 = (~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))) ;
assign n850 = (~((~(n842))*(((~(((n84)*(n208))*(~(n766))))*(~((~(n740))*((n84)*(n208)))))*(~((~(n740))*(~(n766)))))))*(~((n842)*(~(((~(((n84)*(n208))*(~(n766))))*(~((~(n740))*((n84)*(n208)))))*(~((~(n740))*(~(n766)))))))) ;
assign n857 = (~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850))) ;
assign n863 = (~((n690)*((n690)*(~(n850)))))*(~((~(n690))*((~(n690))*(~((~((~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))*(~((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850)))))))*(~((((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850))))))))))) ;
assign n869 = (~((n675)*((n675)*(~(n850)))))*(~((~(n675))*((~(n675))*(~((~((~(((~((n690)*((n690)*(~(n772)))))*(~((~(n690))*((~(n690))*(~((~((~((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782))))))*(~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))))*(~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))))))))*(((~((n690)*((~(n687))*(n690))))*(~((~(n690))*((~(n687))*(~(n690))))))*((~((n690)*((n690)*(~(n782)))))*(~((~(n690))*((~(n690))*(~((~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*(~((n687)*(~((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))))))))))))*(~((~((n690)*((n690)*(~(n850)))))*(~((~(n690))*((~(n690))*(~((~((~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))*(~((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850)))))))*(~((((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850)))))))))))))))*(~((((~((n690)*((n690)*(~(n772)))))*(~((~(n690))*((~(n690))*(~((~((~((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782))))))*(~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))))*(~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))))))))*(((~((n690)*((~(n687))*(n690))))*(~((~(n690))*((~(n687))*(~(n690))))))*((~((n690)*((n690)*(~(n782)))))*(~((~(n690))*((~(n690))*(~((~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*(~((n687)*(~((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))))))))))*((~((n690)*((n690)*(~(n850)))))*(~((~(n690))*((~(n690))*(~((~((~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))*(~((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850)))))))*(~((((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*((~((~((n772)*((n687)*(n782))))*(~(n850))))*(~(((n772)*((n687)*(n782)))*(n850))))))))))))))))))) ;
assign n874 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n97)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n109))) ;
assign n3242 = (((~((~(n16))*((n537)*(~(n540)))))*((~(n557))*(~((n513)*(n534)))))*(~((n513)*(n534))))*(n534) ;
assign n883 = (~((((~((~(n593))*(~(n661))))*(n661))*(~(n874)))*(n3242)))*(~((((~(n593))*(~(n661)))*(n1))*(~(n661)))) ;
assign n898 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n95)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n107))) ;
assign n3252 = (((~((~(n16))*((n537)*(~(n540)))))*((~(n557))*(~((n513)*(n534)))))*(~((n513)*(n534))))*(n534) ;
assign n907 = (~((((~((~(n593))*(~(n661))))*(n661))*(~(n898)))*(n3252)))*(~((((~(n593))*(~(n661)))*(n3))*(~(n661)))) ;
assign n912 = ((~((~((~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208)))))))))))))*(n713)))*(~(((~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208))))))))))))*(~(n713)))))*(~(n673)) ;
assign n3259 = ((~((~((~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))))))*(~((~((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208)))))))))*(~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))))))))))))))*(n907)))*(~(((~(((~(n84))*(n208))*(((~(n84))*(n208))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((~(n84))*(n208)))*((~((~(n84))*(n208)))*(~((~(((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208))))))))*((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734)))))))))))))))))))))))*(~((~((~(((n84)*(~(n208)))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((n84)*(~(n208))))))*(~((~((n84)*(~(n208))))*((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((n84)*(~(n208)))))))))*(~((~(((n84)*(~(n208)))*(((n84)*(~(n208)))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))*(~((~((n84)*(~(n208))))*((~((n84)*(~(n208))))*(~((~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))*(~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*(~((~(((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))))*((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))*(~((~((~(((~(n84))*(n208))*((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*(~((~((~(n84))*(n208)))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))))*(~((~((~(((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))))*(~((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))*(~((((~(n84))*(n208))*(~((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))))*((~(((n84)*(~(n208)))*(n734)))*(~((~((n84)*(~(n208))))*(~(n734))))))))))))))))))))))))))))))*(~(n907)))))*(~((~(n84))*(~(n208)))) ;
assign n916 = (((((~((~(n809))*(n823)))*(~((n809)*(~(n823)))))*(~((~(n869))*(n883))))*(~((n869)*(~(n883)))))*(n3259))*(n912) ;
assign n946 = (~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))) ;
assign n960 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~((~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))*(~(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))))*(~(((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))*(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))))))) ;
assign n970 = (~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))) ;
assign n976 = (~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~((((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))) ;
assign n982 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))*(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))*(~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~((((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))*(~((((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))*(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~(((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))*(~((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))*(~((((~((~((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*((~((~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))))))))*(~(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))*(~(((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(~(((~(((n83)*(n209))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((n83)*(n209)))))*(~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~((~(((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))*((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))*(~((((~(((n83)*(~(n209)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))*(~(((n83)*(~(n209)))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~(((n83)*(n209))*((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))*(~((~((n83)*(n209)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))))))*(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))))))) ;
assign n992 = (~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*(~((~(((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209))))))))*((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))))))))))))))))))*(~((~((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((n83)*(~(n209)))))))))*(~((~(((n83)*(~(n209)))*(((n83)*(~(n209)))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))*(~((~((n83)*(~(n209))))*((~((n83)*(~(n209))))*(~((~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))*(~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~(((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))*(~((~((~(((~(n83))*(n209))*((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))*(~((~((~(n83))*(n209)))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~((~((~((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))*(~(((~(((n83)*(~(n209)))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((n83)*(~(n209))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(((~(n83))*(n209))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))))))))))))))))))))))))))) ;
assign n3266 = (((((~((n823)*(~(n960))))*(~((~(n823))*(n960))))*(~((n883)*(~(n982)))))*(~((~(n883))*(n982))))*(~((n907)*(~(n992)))))*(~((~(n907))*(n992))) ;
assign n1001 = ((((~((n713)*(~((~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681)))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))*(~((n83)*(~(n209)))))))))))))))*(~((~(n713))*((~(((~(n83))*(n209))*(((~(n83))*(n209))*(~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681)))))))))*(~((~((~(n83))*(n209)))*((~((~(n83))*(n209)))*((~(((n83)*(~(n209)))*((~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))*((n83)*(~(n209))))))*(~((~((n83)*(~(n209))))*((~((~(((~(n83))*(n209))*(n681)))*(~((~((~(n83))*(n209)))*(~(n681))))))*(~((n83)*(~(n209)))))))))))))))*(~(n673)))*(~((~(n83))*(~(n209)))))*(n3266) ;
assign n1022 = (~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))) ;
assign n1055 = (~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))) ;
assign n3276 = (((~((n823)*(~((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*(~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))*(~(((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))))))))))*(~((~(n823))*((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))*(~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))*(~(((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))))))))))*(~((n883)*(~((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((~(((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))))))))))*(~((~(n883))*((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~((~(((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))*(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))))))))) ;
assign n3275 = (((~((n713)*(~((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))))))))*(~((~(n713))*((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))))))))*(~(n673)))*(~((~(n82))*(~(n210)))) ;
assign n3274 = ((~((n907)*(~((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))))))))))*(~((~(n907))*((~(((~(n82))*(n210))*(((~(n82))*(n210))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((~(n82))*(n210)))*((~((~(n82))*(n210)))*(~((~(((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210))))))))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))*(~((~((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))))))))))*(n3275) ;
assign n1086 = (n3274)*(n3276) ;
assign n3282 = ((((~((~(n11))*(~(n12))))*(~(n673)))*(n713))*(n823))*(n883) ;
assign n3289 = (((((n11)*(n12))*(~(n673)))*(n713))*(n823))*(n883) ;
assign n3291 = (((((n82)*(n210))*(~((n823)*(~(n1022)))))*(~((~(n823))*(n1022))))*(~((n883)*(~(n1055)))))*(~((~(n883))*(n1055))) ;
assign n1114 = (((~((n907)*(~((~((n681)*(n727)))*(~((~(n681))*(~(n727))))))))*(~((~(n907))*((~((n681)*(n727)))*(~((~(n681))*(~(n727))))))))*(((~((n681)*(n713)))*(~((~(n681))*(~(n713)))))*(~(n673))))*(n3291) ;
assign n3298 = ((((~((n823)*(~((~((~(n766))*(~((n684)*(n734)))))*(~((n766)*((n684)*(n734))))))))*(~((~(n823))*((~((~(n766))*(~((n684)*(n734)))))*(~((n766)*((n684)*(n734))))))))*(~((n907)*(~((~((n684)*(n734)))*(~((~(n684))*(~(n734)))))))))*(~((~(n907))*((~((n684)*(n734)))*(~((~(n684))*(~(n734))))))))*(n747) ;
assign n1131 = (((((~((n684)*(n713)))*(~((~(n684))*(~(n713)))))*(~(n673)))*(~((n883)*(~(n970)))))*(~((~(n883))*(n970))))*(n3298) ;
assign n3305 = ((((~((~((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782))))))*(n823)))*(~(((~((~(n772))*(~((n687)*(n782)))))*(~((n772)*((n687)*(n782)))))*(~(n823)))))*(~((~((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))*(n907))))*(~(((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))*(~(n907)))))*(n741) ;
assign n1148 = (((((~((n687)*(n713)))*(~((~(n687))*(~(n713)))))*(~(n673)))*(~((~(n857))*(n883))))*(~((n857)*(~(n883)))))*(n3305) ;
assign n3314 = ((((n534)*(~(n673)))*(~(n916)))*(~((n907)*(n3282))))*(~((~(n907))*(n3289))) ;
assign n3325 = ((~((~((~((n690)*((n690)*(~(n782)))))*(~((~(n690))*((~(n690))*(~((~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*(~((n687)*(~((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))))))))))*(n907)))*(~(((~((n690)*((n690)*(~(n782)))))*(~((~(n690))*((~(n690))*(~((~((~(n687))*((~((n687)*(n782)))*(~((~(n687))*(~(n782)))))))*(~((n687)*(~((~((n687)*(n782)))*(~((~(n687))*(~(n782))))))))))))))*(~(n907)))))*(((~((~((~((n690)*((~(n687))*(n690))))*(~((~(n690))*((~(n687))*(~(n690)))))))*(n713)))*(~(((~((n690)*((~(n687))*(n690))))*(~((~(n690))*((~(n687))*(~(n690))))))*(~(n713)))))*(~(n673))) ;
assign n1173 = (((((~((~(n795))*(n823)))*(~((n795)*(~(n823)))))*(~((~(n863))*(n883))))*(~((n863)*(~(n883)))))*(n84))*(n3325) ;
assign n3330 = ((~((n907)*(~((~((n717)*((n717)*(~(n734)))))*(~((~(n717))*((~(n717))*(~((~((~(n684))*((~((n684)*(n734)))*(~((~(n684))*(~(n734)))))))*(~((n684)*(~((~((n684)*(n734)))*(~((~(n684))*(~(n734)))))))))))))))))*(~((~(n907))*((~((n717)*((n717)*(~(n734)))))*(~((~(n717))*((~(n717))*(~((~((~(n684))*((~((n684)*(n734)))*(~((~(n684))*(~(n734)))))))*(~((n684)*(~((~((n684)*(n734)))*(~((~(n684))*(~(n734)))))))))))))))))*(((~((n713)*(~((~((n717)*((~(n684))*(n717))))*(~((~(n717))*((~(n684))*(~(n717)))))))))*(~((~(n713))*((~((n717)*((~(n684))*(n717))))*(~((~(n717))*((~(n684))*(~(n717)))))))))*(~(n673))) ;
assign n1190 = (((((~((n823)*(~(n946))))*(~((~(n823))*(n946))))*(~((n883)*(~(n976)))))*(~((~(n883))*(n976))))*(n83))*(n3330) ;
assign n3338 = (((~((n823)*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((~(n823))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((n883)*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))))))))))))*(~((~(n883))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~(((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))))*(~((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))*(~((((~((~((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12)))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*((~((~((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12)))))))))))*(~(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))))))*(~(((~(((~(n11))*(~(n12)))*(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))*(~((~((~(n11))*(~(n12))))*(~(((~(((n82)*(n210))*((~(n11))*(~(n12)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((n82)*(n210)))))*(~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(n11))*(~(n12))))))))))*(((~((~(((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12))))))))*((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))*(~((((~(((n82)*(~(n210)))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))*(~(((n82)*(~(n210)))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~((~(((n82)*(n210))*(~((~(n11))*(~(n12))))))*(~((~((n82)*(n210)))*((~(n11))*(~(n12))))))))))*(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))) ;
assign n3337 = (((~((n713)*(~((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))))*(~((~(n713))*((~(((n82)*(~(n210)))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((n82)*(~(n210))))))*(~((~((n82)*(~(n210))))*((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((n82)*(~(n210)))))))))))*(~(n673)))*(n82) ;
assign n3336 = ((~((n907)*(~((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(~((~(n907))*((~(((n82)*(~(n210)))*(((n82)*(~(n210)))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))*(~((~((n82)*(~(n210))))*((~((n82)*(~(n210))))*(~((~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))*(~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*(~((~(((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12))))))*((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))*(~((~((~(((~(n82))*(n210))*((~(n11))*(n12))))*(~((~((~(n82))*(n210)))*(~((~(n11))*(n12)))))))*(~((~((~((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12)))))))))*(~(((~(n82))*(n210))*(~((~(n11))*(n12)))))))*(~(((~(((n82)*(~(n210)))*(~((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(~((~((n82)*(~(n210))))*((~((~(n11))*(n12)))*(~((n11)*(~(n12))))))))*(((~(n82))*(n210))*(~((~(n11))*(n12)))))))))))))))))))))))*(n3337) ;
assign n1207 = (n3336)*(n3338) ;
assign n1212 = (((((n11)*(~(n673)))*(~(n713)))*(n823))*(n883))*(n907) ;
assign n3351 = (((((n11)*(n12))*(~(n673)))*(~(n713)))*(n823))*(n883) ;
assign n3352 = (((((~((~(n760))*(n823)))*(~((n760)*(~(n823)))))*(~((~(n834))*(n883))))*(~((n834)*(~(n883)))))*(~((~(n727))*(n907))))*(~((n727)*(~(n907)))) ;
assign n1235 = ((((~((~(n681))*(n713)))*(~((n681)*(~(n713)))))*(~(n673)))*((n82)*(n210)))*(n3352) ;
assign n3358 = ((((~((~((~((n676)*(n681)))*(~((~(n676))*(~(n681))))))*(n713)))*(~(((~((n676)*(n681)))*(~((~(n676))*(~(n681)))))*(~(n713)))))*(~(n673)))*(~((~(n766))*(n823))))*(~((n766)*(~(n823)))) ;
assign n1252 = (((((~((~(n842))*(n883)))*(~((n842)*(~(n883)))))*(~((~(n734))*(n907))))*(~((n734)*(~(n907)))))*(n747))*(n3358) ;
assign n3367 = (((((~((~(n687))*(n713)))*(~((n687)*(~(n713)))))*(~(n673)))*(~((~(n772))*(n823))))*(~((n772)*(~(n823)))))*(n741) ;
assign n1269 = ((((~((~(n850))*(n883)))*(~((n850)*(~(n883)))))*(~((~(n782))*(n907))))*(~((n782)*(~(n907)))))*(n3367) ;
assign n3372 = ((~((n3336)*(n3338)))*(~((~(n907))*(n3351))))*((n534)*(~(n1173))) ;
assign n3381 = ((~((~((~(n8))*(n167)))*((n31)*(n53))))*((~((n53)*(n163)))*(~((n53)*(n72)))))*(~((n31)*(n53))) ;
assign n3380 = ((~(((~(((~(n8))*(n44))*(n182)))*(n53))*(n75)))*(~((n53)*(n75))))*(~((n53)*(n150))) ;
assign n1304 = (((n10)*(~(n59)))*(n60))*(n65) ;
assign n1307 = (n34)*(n35) ;
assign n1309 = (n37)*((n36)*((n34)*(n35))) ;
assign n1311 = ((n59)*(~(n60)))*(n65) ;
assign n1313 = ((~(((n59)*(~(n60)))*(n65)))*(~(n178)))*(n200) ;
assign n1321 = ((((~((n907)*(n3282)))*(~((~(n907))*(n3289))))*(~((~(n907))*(n3351))))*(n534))*(~(n1212)) ;
assign n1329 = (n747)*(~(((((n534)*(~(n1001)))*(~(n1131)))*(~(n1190)))*(~(n1252)))) ;
assign n1334 = (((((~(n193))*(n533))*(~(n916)))*(~(n1148)))*(~(n1173)))*(~(n1269)) ;
assign n3403 = (((~((n3274)*(n3276)))*(~((n3336)*(n3338))))*(n534))*(~(n1114)) ;
assign n3404 = (~(((n11)*(n12))*(~(n1321))))*(~(((n84)*(n208))*(~(n1334)))) ;
assign n1344 = ((~(((n82)*(n210))*(~((~(n1235))*(n3403)))))*(~(n1329)))*(n3404) ;
assign n3412 = (~((~(((~((~(n487))*(~(n544))))*(n111))*(n567)))*(~((((~(n487))*(~(n544)))*(n121))*(~(n567))))))*(n534) ;
assign n1358 = (~((((~(n542))*(~(n557)))*(~(n578)))*(n3412)))*(~(((n137)*(n578))*(n583))) ;
assign n1363 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1358))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n140))*(~(n661)))) ;
assign n3420 = (~((~(((~((~(n487))*(~(n544))))*(n112))*(n567)))*(~((((~(n487))*(~(n544)))*(n122))*(~(n567))))))*(n534) ;
assign n1377 = (~((((~(n542))*(~(n557)))*(~(n578)))*(n3420)))*(~(((n138)*(n578))*(n583))) ;
assign n1382 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1377))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n141))*(~(n661)))) ;
assign n3428 = (~((~(((~((~(n487))*(~(n544))))*(n110))*(n567)))*(~((((~(n487))*(~(n544)))*(n120))*(~(n567))))))*(n534) ;
assign n1396 = (~((((~(n542))*(~(n557)))*(~(n578)))*(n3428)))*(~(((n136)*(n578))*(n583))) ;
assign n1401 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1396))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n139))*(~(n661)))) ;
assign n1406 = (((((~(n13))*(n1313))*(~(n1363)))*(~(n1382)))*(~(n1401)))*(~(n1344)) ;
assign n1407 = (n120)*(n122) ;
assign n1408 = (n124)*((n120)*(n122)) ;
assign n3438 = (((n126)*((n124)*((n120)*(n122))))*(n121))*(n123) ;
assign n1414 = (((n125)*(n127))*(n128))*(n3438) ;
assign n1420 = (~((~(n70))*(~(n77))))*(~((~(n513))*(~((n58)*(~(n545)))))) ;
assign n1421 = (~((n169)*(~((n168)*((~(n17))*(n485))))))*(~((~(n549))*((~(n537))*(~((~(n17))*(n485)))))) ;
assign n1426 = (n30)*(((((~(n54))*(~(n55)))*(n56))*(n29))*(~(n57))) ;
assign n1429 = (~((n67)*((n66)*((((n29)*(~(n30)))*(~(n57)))*(n599)))))*(~((~(n67))*((~(n66))*((((~(n57))*(n599))*(~(n29)))*(~(n30)))))) ;
assign n1431 = (~((n30)*(((n29)*(~(n57)))*(n544))))*(~((~(n627))*(~(n1429)))) ;
assign n1435 = (n5)*(~((((~((~(n626))*(n627)))*(~((n627)*(n630))))*(~(n17)))*(n1431))) ;
assign n3447 = ((((~((n30)*(((~(n29))*(~(n57)))*(n544))))*(~((~(n30))*(((~(n29))*(~(n57)))*(n544)))))*(~((~(n30))*(((n29)*(~(n57)))*(n544)))))*((~((n57)*(n544)))*(n626)))*(~((n57)*(n599))) ;
assign n1443 = ((~(((n58)*(~((~(n487))*(~(n544)))))*(~(n1429))))*(~((~(n626))*(~((n58)*(~((~(n487))*(~(n544)))))))))*(n647) ;
assign n3451 = ((~((~(n501))*(~((n534)*(n3447)))))*(~((n16)*(~((n534)*(n1443))))))*(~((n20)*(~(n534)))) ;
assign n3450 = (~((((~(n18))*(n19))*(n513))*(~(n1311))))*(~((~(n501))*(n1421))) ;
assign n1454 = ((((~((n15)*(n628)))*(~(n1313)))*(~(n1435)))*(n3450))*(n3451) ;
assign n1457 = (~(n64))*(((n59)*(~(n60)))*(n65)) ;
assign n3466 = ((~((((~(n13))*(n38))*(n1309))*(n1313)))*(~((n1313)*(n1457))))*(~((n40)*(n1313))) ;
assign n3465 = (((~((n1454)*(~((n13)*(n1313)))))*(~(n22)))*(~(n1420)))*(~(((~(n13))*(n1313))*(n1414))) ;
assign n3474 = (~((n16)*(~(((~((n627)*(~(n1429))))*(~((~(n626))*(~(n627)))))*(n647)))))*(~((n15)*((~(n626))*(n627)))) ;
assign n1476 = (~((~(n204))*(n205)))*(~((n204)*(n205))) ;
assign n3479 = (((~((~(n3))*(~((~((~((n675)*(~(n684))))*(~((~((n690)*(n734)))*(~((~(n690))*(~(n734))))))))*(~(((n675)*(~(n684)))*((~((n690)*(n734)))*(~((~(n690))*(~(n734)))))))))))*(~((n3)*((~((~((n675)*(~(n684))))*(~((~((n690)*(n734)))*(~((~(n690))*(~(n734))))))))*(~(((n675)*(~(n684)))*((~((n690)*(n734)))*(~((~(n690))*(~(n734)))))))))))*((~((n675)*(n684)))*(~((~(n675))*(~(n684))))))*(n4) ;
assign n3486 = ((~(((((~((~(n1))*(~(n850))))*(~((n1)*(n850))))*((~((~(n2))*(~(n772))))*(~((n2)*(n772)))))*(n3))*(n782)))*(~((((~((~(n1))*(~(n850))))*(~((n1)*(n850))))*(n2))*(n772))))*(~((n1)*(n850))) ;
assign n1500 = (~((((~((~(n1))*(~(n850))))*(~((n1)*(n850))))*((~((~(n2))*(~(n772))))*(~((n2)*(n772)))))*(n3479)))*(n3486) ;
assign n1504 = (n19)*((n28)*((~(n30))*(n596))) ;
assign n1510 = (~(n30))*((((~(n27))*(n29))*(~(n57)))*(n489)) ;
assign n1511 = (n28)*((~(n30))*((((~(n27))*(n29))*(~(n57)))*(n489))) ;
assign n1513 = (n28)*((~(n30))*((((n27)*(n29))*(~(n57)))*(n489))) ;
assign n1514 = (~(n28))*((~(n30))*((((n27)*(n29))*(~(n57)))*(n489))) ;
assign n1518 = (n5)*(~((((~((~(n17))*((n28)*((n30)*(n492)))))*(~((n28)*((~(n30))*(n497)))))*(~((n28)*((~(n30))*(n492)))))*(~((~(n28))*((~(n30))*(n492)))))) ;
assign n3495 = ((~(((~((~(n538))*(~(n599))))*(~(n501)))*(~(n513))))*(~((n19)*(n513))))*(~((~(n501))*(n544))) ;
assign n1523 = (~(n1500))*(~(((~(n1504))*(~(n1518)))*(n3495))) ;
assign n1541 = (~((~((~((n141)*(~(n142))))*(~((~(n141))*(n142)))))*((~((n143)*(~(n144))))*(~((~(n143))*(n144))))))*(~(((~((n141)*(~(n142))))*(~((~(n141))*(n142))))*(~((~((n143)*(~(n144))))*(~((~(n143))*(n144))))))) ;
assign n1547 = (~((n257)*((~((~((~((~((~((~(n66))*(n67)))*(~((n66)*(~(n67))))))*((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))*(~(((~((~(n66))*(n67)))*(~((n66)*(~(n67)))))*(~((~((n139)*(~(n140))))*(~((~(n139))*(n140)))))))))*(n1541)))*(~(((~((~((~((~(n66))*(n67)))*(~((n66)*(~(n67))))))*((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))*(~(((~((~(n66))*(n67)))*(~((n66)*(~(n67)))))*(~((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))))*(~(n1541)))))))*(~((~(n257))*(~((~((~((~((~((~((~(n66))*(n67)))*(~((n66)*(~(n67))))))*((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))*(~(((~((~(n66))*(n67)))*(~((n66)*(~(n67)))))*(~((~((n139)*(~(n140))))*(~((~(n139))*(n140)))))))))*(n1541)))*(~(((~((~((~((~(n66))*(n67)))*(~((n66)*(~(n67))))))*((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))*(~(((~((~(n66))*(n67)))*(~((n66)*(~(n67)))))*(~((~((n139)*(~(n140))))*(~((~(n139))*(n140))))))))*(~(n1541)))))))) ;
assign n1565 = (~((~((~((~(n247))*(n248)))*(~((n247)*(~(n248))))))*((~((n254)*(~(n255))))*(~((~(n254))*(n255))))))*(~(((~((~(n247))*(n248)))*(~((n247)*(~(n248)))))*(~((~((n254)*(~(n255))))*(~((~(n254))*(n255))))))) ;
assign n1571 = (~((n256)*((~((~((~((~((~((n145)*(~(n146))))*(~((~(n145))*(n146)))))*((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))*(~(((~((n145)*(~(n146))))*(~((~(n145))*(n146))))*(~((~((n147)*(~(n148))))*(~((~(n147))*(n148)))))))))*(n1565)))*(~(((~((~((~((n145)*(~(n146))))*(~((~(n145))*(n146)))))*((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))*(~(((~((n145)*(~(n146))))*(~((~(n145))*(n146))))*(~((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))))*(~(n1565)))))))*(~((~(n256))*(~((~((~((~((~((~((n145)*(~(n146))))*(~((~(n145))*(n146)))))*((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))*(~(((~((n145)*(~(n146))))*(~((~(n145))*(n146))))*(~((~((n147)*(~(n148))))*(~((~(n147))*(n148)))))))))*(n1565)))*(~(((~((~((~((n145)*(~(n146))))*(~((~(n145))*(n146)))))*((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))*(~(((~((n145)*(~(n146))))*(~((~(n145))*(n146))))*(~((~((n147)*(~(n148))))*(~((~(n147))*(n148))))))))*(~(n1565)))))))) ;
assign n1576 = (n28)*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489))) ;
assign n1579 = (n5)*(~(((~(n598))*(~(n1514)))*(~(n1576)))) ;
assign n1580 = (~(((~(n54))*(~(n55)))*(n56)))*(~((~(n17))*(((~(n54))*(~(n55)))*(~(n56))))) ;
assign n1584 = (~((~(n1547))*(~(n1571))))*(~((~(n1579))*(~((~(n501))*(~((~(n538))*(n1580))))))) ;
assign n1586 = (n188)*(~((n5)*(n178))) ;
assign n3501 = (((~((n18)*(n19)))*((~(n21))*(~(n22))))*(n534))*(~(n1420)) ;
assign n3510 = ((~((((~(n13))*(n38))*(n1309))*(n1313)))*(~(((~(n13))*(n1313))*(n1414))))*(~((n1313)*(n1457))) ;
assign n3509 = (((((n1476)*(~(n1523)))*(~(n1584)))*(~(n1586)))*(n3501))*(~(n1406)) ;
assign n1601 = ((((~((n40)*(n1313)))*(~((n1304)*(n1313))))*(~(n1454)))*(n3509))*(n3510) ;
assign n1604 = (~(n549))*(~((n202)*(~((~(n537))*(~((~(n17))*(n485))))))) ;
assign n1608 = ((~((~(n17))*(((((n30)*(~(n54)))*(n55))*(n56))*(~(n57)))))*(~(((((~(n30))*(~(n54)))*(n55))*(n56))*(~(n57)))))*(~((((~(n54))*(n55))*(n56))*(n57))) ;
assign n3523 = (~((~((~(n70))*(~(n77))))*((n540)*(~(n1608)))))*(~(((n16)*(n540))*(~(n1604)))) ;
assign n1616 = ((~(((~((n5)*(n598)))*(~(n41)))*(n3523)))*(~((n15)*(n598))))*(~(n40)) ;
assign n1620 = ((~(n28))*((~(n30))*(n492)))*(~(n1584)) ;
assign n1621 = (~((n58)*(~((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(~(n55)))*(n56)))))))*((n57)*((~(n17))*(((~(n54))*(~(n55)))*(~(n56))))) ;
assign n1626 = (n5)*(~(((((~(n537))*(~(n538)))*(~(n591)))*(~(n1620)))*(~(n1621)))) ;
assign n1628 = (~((n28)*((~(n30))*((((~(n27))*(n29))*(~(n57)))*(n489)))))*(~((n28)*((~(n30))*((((n27)*(n29))*(~(n57)))*(n489))))) ;
assign n3535 = ((~((n5)*(~((~(n1511))*(~(n1513))))))*(~((n16)*(n631))))*(~((n15)*(n1513))) ;
assign n3540 = (((~((n15)*((~(n626))*(n627))))*(~(((n16)*(~(n626)))*(~(n627)))))*(~((n5)*((~(n627))*(~(n1429))))))*(~((n16)*((n627)*(~(n1429))))) ;
assign n3539 = (~((n5)*((n30)*(((n29)*(~(n57)))*(n544)))))*(~((n16)*(~(((~((n30)*(((~(n29))*(~(n57)))*(n544))))*(~((~(n30))*(((~(n29))*(~(n57)))*(n544)))))*(~((~(n30))*(((n29)*(~(n57)))*(n544)))))))) ;
assign n1668 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n93)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n105))) ;
assign n1672 = (~((((~((~(n193))*(n533)))*(n52))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1668)))) ;
assign n1679 = (~((((~((n513)*(n534)))*(~((~(n593))*(~(n661)))))*(n661))*(~(n1672))))*(~((((~(n593))*(~(n661)))*(n135))*(~(n661)))) ;
assign n1688 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n92)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n104))) ;
assign n1692 = (~((((~((~(n193))*(n533)))*(n130))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1688)))) ;
assign n1702 = (~(((~((~((~(n578))*((~(n578))*(~(n1692)))))*(~((n578)*((n578)*(~(n583)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n134))*(~(n661)))) ;
assign n1711 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n91)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n103))) ;
assign n1715 = (~((((~((~(n193))*(n533)))*(n49))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1711)))) ;
assign n1725 = (~(((~((~((~(n578))*((~(n578))*(~(n1715)))))*(~((n578)*((n578)*(n583))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n133))*(~(n661)))) ;
assign n1734 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n90)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n102))) ;
assign n1738 = (~((((~((~(n193))*(n533)))*(n50))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1734)))) ;
assign n1745 = ((n513)*(n534))*(((n513)*(n534))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n1)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))))))) ;
assign n1751 = (~(((~((~((~(n578))*((~(n578))*(~(n1738)))))*(~(n1745))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n132))*(~(n661)))) ;
assign n1760 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n89)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n101))) ;
assign n1764 = (~((((~((~(n193))*(n533)))*(n48))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1760)))) ;
assign n1771 = ((n513)*(n534))*(((n513)*(n534))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n2)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))))))) ;
assign n1777 = (~(((~((~((~(n578))*((~(n578))*(~(n1764)))))*(~(n1771))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n131))*(~(n661)))) ;
assign n1786 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n88)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n100))) ;
assign n1790 = (~((((~((~(n193))*(n533)))*(n51))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1786)))) ;
assign n1797 = ((n513)*(n534))*(((n513)*(n534))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n3)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))))))) ;
assign n1803 = (~(((~((~((~(n578))*((~(n578))*(~(n1790)))))*(~(n1797))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n138))*(~(n661)))) ;
assign n1812 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n87)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n99))) ;
assign n1816 = (~((((~((~(n193))*(n533)))*(n47))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1812)))) ;
assign n1822 = (~((n1)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n4)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n1830 = (~(((~((~((~(n578))*((~(n578))*(~(n1816)))))*(~((n578)*((n578)*(~(n1822)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n137))*(~(n661)))) ;
assign n1836 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n86)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n98))) ;
assign n1840 = (~((((~((~(n193))*(n533)))*(n52))*(~(n542)))*(n557)))*(~(((((~(n193))*(n533))*(~(n542)))*(~(n557)))*(~(n1836)))) ;
assign n1846 = (~((n2)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n135)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n1854 = (~(((~((~((~(n578))*((~(n578))*(~(n1840)))))*(~((n578)*((n578)*(~(n1846)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n136))*(~(n661)))) ;
assign n1858 = (n129)*((((n125)*(n127))*(n128))*(n3438)) ;
assign n1860 = ((~((n28)*((n30)*(n596))))*(n24))*(~(n43)) ;
assign n1864 = ((((n244)*(n245))*(n540))*(~(n1858)))*(n1860) ;
assign n1865 = (~(((n501)*(~(n540)))*(~(n567))))*(~(n1864)) ;
assign n3631 = ((~((~(n501))*((~(n17))*(n485))))*(~((~(n501))*(n537))))*(~((~((~(n120))*(n121)))*(~((n120)*(~(n121)))))) ;
assign n3638 = ((~((~((n122)*(~((n120)*(n121)))))*(~((~(n122))*((n120)*(n121))))))*(~((~(n501))*(n537))))*(~((~(n501))*(n538))) ;
assign n1903 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n113)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n123))) ;
assign n1912 = (~((n131)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n136)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n1915 = (~(((((~((n513)*(n534)))*(n534))*(~(n542)))*(~(n557)))*(~(n1903))))*(~(((n513)*(n534))*(((n513)*(n534))*(~(n1912))))) ;
assign n1920 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1915))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n142))*(~(n661)))) ;
assign n3650 = (~((~((n123)*(~((n121)*((n120)*(n122))))))*(~((~(n123))*((n121)*((n120)*(n122)))))))*(~((~(n501))*(n537))) ;
assign n1937 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n114)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n124))) ;
assign n1946 = (~((n132)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n137)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n1949 = (~(((((~((n513)*(n534)))*(n534))*(~(n542)))*(~(n557)))*(~(n1937))))*(~(((n513)*(n534))*(((n513)*(n534))*(~(n1946))))) ;
assign n1954 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1949))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n143))*(~(n661)))) ;
assign n3666 = (~((~((n124)*(~((((n120)*(n122))*(n121))*(n123)))))*(~((~(n124))*((((n120)*(n122))*(n121))*(n123))))))*(~(n1865)) ;
assign n1972 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n115)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n125))) ;
assign n1981 = (~((n133)*((n513)*(~(((~(n5))*(~(n16)))*(~(n164)))))))*(~((~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))*((n138)*(~((n513)*(~(((~(n5))*(~(n16)))*(~(n164))))))))) ;
assign n1984 = (~(((((~((n513)*(n534)))*(n534))*(~(n542)))*(~(n557)))*(~(n1972))))*(~(((n513)*(n534))*(((n513)*(n534))*(~(n1981))))) ;
assign n1989 = (~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1984))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n144))*(~(n661)))) ;
assign n1998 = (~((n125)*(~((((n124)*((n120)*(n122)))*(n121))*(n123)))))*(~((~(n125))*((((n124)*((n120)*(n122)))*(n121))*(n123)))) ;
assign n2012 = (~((n126)*(~(((((n124)*(n1407))*(n121))*(n123))*(n125)))))*(~((~(n126))*(((((n124)*(n1407))*(n121))*(n123))*(n125)))) ;
assign n2020 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n116)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n126))) ;
assign n3694 = (((~((n169)*(~((n168)*(n538)))))*(~(n16)))*(n27))*(n534) ;
assign n2029 = (~((((n534)*(~(n542)))*(~(n557)))*(~(n2020))))*(~(((n537)*(n557))*(n3694))) ;
assign n2038 = (~((~((n513)*(n534)))*((~((n513)*(n534)))*(~(n2029)))))*(~(((n513)*(n534))*(((n513)*(n534))*(~((~((n134)*(n583)))*(~((~(n583))*((n131)*(~(n583)))))))))) ;
assign n2043 = (~(((~((~(n593))*(~(n661))))*(n661))*(~(n2038))))*(~((((~(n593))*(~(n661)))*(n145))*(~(n661)))) ;
assign n3701 = (~(((((~((~(n501))*(n538)))*(n27))*(~(n501)))*(n537))*(n1865)))*(~((((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(~(n1865)))*(~(n2012)))) ;
assign n2059 = (~((n127)*(~(((((n126)*(n1408))*(n121))*(n123))*(n125)))))*(~((~(n127))*(((((n126)*(n1408))*(n121))*(n123))*(n125)))) ;
assign n2067 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n117)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n127))) ;
assign n3718 = (((~((n169)*(~((n168)*(n538)))))*(~(n16)))*(n28))*(n534) ;
assign n2076 = (~((((n534)*(~(n542)))*(~(n557)))*(~(n2067))))*(~(((n537)*(n557))*(n3718))) ;
assign n2085 = (~((~((n513)*(n534)))*((~((n513)*(n534)))*(~(n2076)))))*(~(((n513)*(n534))*(((n513)*(n534))*(~((~((n135)*(n583)))*(~((~(n583))*((n132)*(~(n583)))))))))) ;
assign n2090 = (~(((~((~(n593))*(~(n661))))*(n661))*(~(n2085))))*(~((((~(n593))*(~(n661)))*(n146))*(~(n661)))) ;
assign n3725 = (~(((((~((~(n501))*(n538)))*(n28))*(~(n501)))*(n537))*(n1865)))*(~((((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(~(n1865)))*(~(n2059)))) ;
assign n3732 = ((((n126)*((n124)*(n1407)))*(n121))*(n123))*(n125) ;
assign n3733 = ((~((~((n128)*(~((n127)*(n3732)))))*(~((~(n128))*((n127)*(n3732))))))*(~((~(n501))*(n537))))*(~((~(n501))*(n538))) ;
assign n2115 = (~(((~((~(n487))*(~(n544))))*((~(n549))*(n566)))*(n118)))*(~((((~(n487))*(~(n544)))*(~((~(n549))*(n566))))*(n128))) ;
assign n3742 = (((~((n169)*(~((n168)*(n538)))))*(~(n16)))*(n29))*(n534) ;
assign n2124 = (~((((n534)*(~(n542)))*(~(n557)))*(~(n2115))))*(~(((n537)*(n557))*(n3742))) ;
assign n2133 = (~((~((n513)*(n534)))*((~((n513)*(n534)))*(~(n2124)))))*(~(((n513)*(n534))*(((n513)*(n534))*(~((~((n4)*(n583)))*(~((~(n583))*((n133)*(~(n583)))))))))) ;
assign n2138 = (~(((~((~(n593))*(~(n661))))*(n661))*(~(n2133))))*(~((((~(n593))*(~(n661)))*(n147))*(~(n661)))) ;
assign n3749 = (~(((((~((~(n501))*(n538)))*(n29))*(~(n501)))*(n537))*(n1865)))*(~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n2138)))) ;
assign n3753 = (~((~((n129)*(~((((n125)*(n127))*(n128))*(n3438)))))*(~((~(n129))*((((n125)*(n127))*(n128))*(n3438))))))*(~(n1865)) ;
assign n3758 = (~(((((~((~(n501))*(n538)))*(n30))*(~(n501)))*(n537))*(n1865)))*(~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(~(n667)))*(n1865))) ;
assign n3775 = (~((((n15)*(~(n22)))*(~(n1311)))*(n1513)))*(~((((~(n22))*(~(n1311)))*(~(n1586)))*(n1626))) ;
assign n2207 = ((((n59)*(~(n60)))*(n65))*(n64))*(~(n79)) ;
assign n2213 = (~(n28))*((~(n30))*((((~(n27))*(n29))*(~(n57)))*(n489))) ;
assign n2216 = ((((~(n28))*(n1510))*(n15))*(~(n544)))*(n1586) ;
assign n2219 = ((((n58)*(~((~(n487))*(~(n544)))))*(n16))*(~(n544)))*(n1586) ;
assign n2221 = ((n18)*(n172))*(n178) ;
assign n3791 = (((~((~(n17))*((n28)*(n493))))*(~((~(n28))*(n1510))))*(~(n544)))*(~(n627)) ;
assign n2225 = ((((~((~(n17))*(n494)))*(~(n544)))*(~(n627)))*(n1586))*(~(n2213)) ;
assign n2228 = ((((~(n17))*(n494))*(n16))*(~(n544)))*(n1586) ;
assign n3799 = ((((~((n1586)*(n3791)))*(~(n22)))*(~(n2216)))*(~(n2219)))*(~(n2221)) ;
assign n2233 = (~(n2228))*(n3799) ;
assign n3802 = (((~((~(n549))*((~(n537))*(~(n538)))))*(~((n5)*(~((~(n537))*(~(n538)))))))*(n201))*(n501) ;
assign n3808 = (((((~(n70))*(~(n77)))*(~(n45)))*(n201))*(n244))*(n245) ;
assign n3810 = (~((((((~(n45))*(n192))*(n246))*(n501))*(n540))*(~(n1604))))*(~((((n192)*(n501))*(~(n540)))*(~(n1604)))) ;
assign n2251 = (((~(((n246)*(n540))*(n3808)))*(~((~(n540))*(n3802))))*(n2233))*(n3810) ;
assign n2254 = (((~(((n64)*(~(n79)))*(n1311)))*(~((~(n64))*(n1311))))*(~(n40)))*(n2251) ;
assign n2259 = (n7)*(~(n8)) ;
assign n2261 = (n5)*(~((~(n494))*(~(n499)))) ;
assign n2263 = (~(n70))*(~((~(n17))*((n5)*(~((~(n494))*(~(n499))))))) ;
assign n2266 = (n32)*((n7)*(~(n8))) ;
assign n2277 = (((((n27)*(~(n29)))*(~(n28)))*(~(n30)))*(n57))*(n489) ;
assign n2278 = (n28)*(((((~(n27))*(~(n29)))*(~(n30)))*(n57))*(n489)) ;
assign n2286 = ((~((((((~(n27))*(~(n28)))*(n29))*(n30))*(~(n57)))*(n489)))*(~(((((~((~(n28))*(((((~(n27))*(~(n29)))*(~(n30)))*(n57))*(n489))))*(~((((((n27)*(~(n29)))*(~(n28)))*(~(n30)))*(n57))*(n489))))*(~((n28)*(((((~(n27))*(~(n29)))*(~(n30)))*(n57))*(n489)))))*(n57))*(n489))))*(~((~(n28))*((~(n30))*((((~(n27))*(~(n29)))*(~(n57)))*(n489))))) ;
assign n2298 = ((~((((~(((n54)*(n55))*(n56)))*(~(((n54)*(~(n55)))*(n56))))*(~(((n54)*(n55))*(~(n56)))))*(n2286)))*(~((~(n40))*(~(n2286)))))*(n534) ;
assign n2301 = (~(n28))*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489))) ;
assign n2306 = (n28)*((~(n30))*((((~(n27))*(~(n29)))*(~(n57)))*(n489))) ;
assign n2307 = (~(n28))*((n30)*((((n27)*(~(n29)))*(~(n57)))*(n489))) ;
assign n2308 = (~(n28))*((~(n30))*((((n27)*(~(n29)))*(~(n57)))*(n489))) ;
assign n3829 = (((((~((n28)*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489)))))*(~((~(n28))*((n30)*((((n27)*(n29))*(~(n57)))*(n489))))))*(~((~(n28))*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489))))))*(~((n28)*((~(n30))*((((~(n27))*(~(n29)))*(~(n57)))*(n489))))))*(~((~(n28))*((n30)*((((n27)*(~(n29)))*(~(n57)))*(n489))))))*(~((~(n28))*((~(n30))*((((n27)*(~(n29)))*(~(n57)))*(n489))))) ;
assign n2314 = (~(((((~(n16))*(n85))*(~(n170)))*(~(n171)))*(~(n534))))*(n3829) ;
assign n2317 = (~((n28)*((~(n30))*((((~(n27))*(n29))*(~(n57)))*(n489)))))*(~((~(n28))*((~(n30))*((((n27)*(n29))*(~(n57)))*(n489))))) ;
assign n2320 = ((~((n5)*(~(n2314))))*(~((n78)*(n1513))))*(~((n15)*(~(n2317)))) ;
assign n2328 = ((((~((~(n1311))*(n2219)))*(~((n79)*(n1311))))*(~((~(n1311))*(n2225))))*(~((~(n1311))*(n2228))))*(~(n2216)) ;
assign n2336 = (~(n22))*(~((~((~(n549))*(~((n202)*(~(n566))))))*(~((~(n1304))*(n2254))))) ;
assign n3837 = (((~(((~((~(n64))*(n1311)))*(~(n2320)))*(n2328)))*(~(((n64)*(~(n79)))*(n1311))))*(~((n79)*(~(n1311)))))*(~(n6)) ;
assign n3851 = ((~((((n5)*(~(n500)))*(n513))*(~(n2263))))*(~((~(n500))*(n509))))*(~((n5)*(~(n2286)))) ;
assign n2366 = (((~((((n5)*(~(n500)))*(n513))*(~(n2263))))*(n5))*(n2286))*(n2314) ;
assign n2369 = (n16)*(~(((~((~(n627))*(n630)))*(n567))*(~(n591)))) ;
assign n2380 = (((((~(n538))*(~(n591)))*(n626))*(~(n630)))*(n647))*(n1429) ;
assign n3868 = ((~((n598)*(~((~(n164))*(~(n181))))))*(~((~(n166))*(n1514))))*(~((n166)*(~(n2380)))) ;
assign n2397 = (n151)*((((~(((n64)*(~(n79)))*(n1311)))*(~((~(n64))*(n1311))))*(~(n40)))*(n2251)) ;
assign n2402 = (((~((~(n17))*(n485)))*(~((~(n627))*(n630))))*(~(n537)))*(~(n1426)) ;
assign n3887 = (((~((~(n17))*(n494)))*(~((~(n17))*(n499))))*((n16)*(~(n1313))))*(n151) ;
assign n3886 = (((~((~(n627))*(~(n1429))))*(~(n549)))*(~(n591)))*(~((~(n28))*(n671))) ;
assign n2413 = (((n2254)*(n2402))*(n3886))*(n3887) ;
assign n3897 = ((~(((~(n17))*(n487))*((n58)*(~((~(n487))*(~(n544)))))))*(~((~(n17))*(n494))))*(~((~(n40))*(n544))) ;
assign n2424 = ((((~((~(n2213))*(n3897)))*(~(n6)))*(n151))*(~(n1311)))*(n1586) ;
assign n3901 = ((~(((((~((~(n2213))*(n3897)))*(~(n6)))*(n151))*(~(n1311)))*(n1586)))*(~(n1311)))*(n1586) ;
assign n2429 = (n485)*((n79)*(((n59)*(~(n60)))*(n65))) ;
assign n2430 = (~(((n485)*(~(n499)))*(n3901)))*(~((n485)*((n79)*(n1311)))) ;
assign n2439 = (~(n1586))*(~(((((~(n61))*(~(n62)))*(~(n63)))*(~(n64)))*(~(n76)))) ;
assign n3911 = ((((~((n627)*(~(n1429))))*(~((~(n626))*(~(n627)))))*(~((n28)*(n1510))))*(~((~(n28))*(n1510))))*(n15) ;
assign n3922 = (((~((((n192)*(n501))*(~(n540)))*(~(n1604))))*(~((n501)*(n1858))))*(~((n501)*(n540))))*(~((n13)*(n501))) ;
assign n3927 = ((((~((((n192)*(n501))*(~(n540)))*(~(n1604))))*(~((n13)*(n501))))*(n501))*(~(n540)))*(n549) ;
assign n2508 = ((~(n5))*(~(n15)))*(~(n180)) ;
assign n2509 = (~((~(n193))*(n533)))*(~(((~(n5))*(~(n15)))*(~(n180)))) ;
assign n3942 = (((((n20)*(~(n61)))*(~(n62)))*(n63))*(n76))*(n513) ;
assign n2535 = (n207)*(((((n158)*(n159))*(n160))*(n161))*(n162)) ;
assign n3956 = (~((((~(n19))*(~(n20)))*(~(n173)))*(~(n174))))*((~(n2228))*(n3799)) ;
assign n3962 = ((~(((n5)*(n179))*(~(n545))))*(~((n5)*(n178))))*(~((n169)*(~(n567)))) ;
assign n3965 = (~((~(n178))*((n5)*(~((~(n1426))*(~((~(n627))*(~(n1429)))))))))*(~((n16)*((n627)*(~(n1429))))) ;
assign n2585 = ((~(((~(n13))*(n177))*(n3962)))*(~((~(n24))*(~(n43)))))*(n3965) ;
assign n2591 = (((~((n544)*(n1586)))*(~(((n5)*(n27))*(n544))))*(n2251))*(~(n2585)) ;
assign n3979 = ((((~((~(n907))*(n3289)))*(~((~(n907))*(n3351))))*(~(n1114)))*(~(n1131)))*(~(n1148)) ;
assign n2603 = ((~((~((n544)*(n1586)))*(~(((n5)*(n27))*(n544)))))*(n2251))*(~(n2261)) ;
assign n3988 = (((~((n3274)*(n3276)))*((~(n1173))*(~(n1269))))*(~(n916)))*(~(n1114)) ;
assign n3997 = (((((~(n1173))*(~(n1269)))*(~(n916)))*(~(n1001)))*(~(n1131)))*(~(n1148)) ;
assign n2657 = (~(((((n230)*(~(n2278)))*(n2301))*(~(n2307)))*((~((((n231)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n217)*(n2278))*(~(n2301)))*(~(n2307)))))))*(~((~((((n230)*(~(n2278)))*(n2301))*(~(n2307))))*(~((~((((n231)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n217)*(n2278))*(~(n2301)))*(~(n2307)))))))) ;
assign n4010 = (~(((((n195)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n153)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n2671 = (~(((((n218)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(n4010) ;
assign n4018 = (~(((((n219)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(~(((((n216)*(n2277))*(~(n2301)))*(~(n2306)))*(~(n2308)))) ;
assign n4017 = (~(((((n196)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n154)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n2690 = (n4017)*(n4018) ;
assign n4024 = (~(((((n220)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(~(((((n215)*(n2277))*(~(n2301)))*(~(n2306)))*(~(n2308)))) ;
assign n4023 = (~(((((n197)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n155)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n4030 = (~(((((n221)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(~(((((n214)*(n2277))*(~(n2301)))*(~(n2306)))*(~(n2308)))) ;
assign n4029 = (~(((((n198)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n156)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n2734 = (n4029)*(n4030) ;
assign n4036 = (~(((((n222)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(~(((((n213)*(n2277))*(~(n2301)))*(~(n2306)))*(~(n2308)))) ;
assign n4035 = (~(((((n199)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n157)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n4042 = (~(((((n223)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(~(((((n212)*(n2277))*(~(n2301)))*(~(n2306)))*(~(n2308)))) ;
assign n4041 = (~(((((n194)*(~(n2277)))*(~(n2301)))*(n2306))*(~(n2308))))*(~(((((n152)*(~(n2277)))*(~(n2301)))*(~(n2306)))*(n2308))) ;
assign n2775 = (n4041)*(n4042) ;
assign n2778 = (~((~((n4035)*(n4036)))*(n2775)))*(~(((n4035)*(n4036))*(~(n2775)))) ;
assign n2781 = (~((~((~((~((n4023)*(n4024)))*(n2734)))*(~(((n4023)*(n4024))*(~(n2734))))))*(n2778)))*(~(((~((~((n4023)*(n4024)))*(n2734)))*(~(((n4023)*(n4024))*(~(n2734)))))*(~(n2778)))) ;
assign n2789 = (~(((n238)*(n1628))*(n2307)))*(~(((n240)*(~(n1628)))*(~(n2307)))) ;
assign n2794 = (~(((n239)*(n1628))*(n2307)))*(~(((n241)*(~(n1628)))*(~(n2307)))) ;
assign n2797 = (~((~(n2789))*(n2794)))*(~((n2789)*(~(n2794)))) ;
assign n2804 = (~((((n224)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n232)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2811 = (~((((n225)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n233)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2824 = (~((((n226)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n234)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2831 = (~((((n227)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n235)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2841 = (~((((n228)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n236)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2848 = (~((((n229)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n237)*(~(n2278)))*(~(n2301)))*(n2307))) ;
assign n2851 = (~((~(n2841))*(n2848)))*(~((n2841)*(~(n2848)))) ;
assign n2867 = (n1514)*(~((~((n15)*(n186)))*(~((n16)*(n185))))) ;
assign n4069 = (~(((n169)*(~((n168)*(n538))))*(~(((~(n537))*(~(n538)))*(~(n549))))))*(~(n6)) ;
assign n2884 = ((~((((~(n16))*(n85))*(~(n170)))*(~(n171))))*(n151))*(n193) ;
assign n4075 = (((((~((n28)*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489)))))*(~((~(n28))*((n30)*((((n27)*(n29))*(~(n57)))*(n489))))))*(~((~(n28))*((n30)*((((~(n27))*(~(n29)))*(~(n57)))*(n489))))))*(~((n28)*((~(n30))*((((~(n27))*(~(n29)))*(~(n57)))*(n489))))))*(~((~(n28))*((n30)*((((n27)*(~(n29)))*(~(n57)))*(n489))))))*(~((~(n28))*((~(n30))*((((n27)*(~(n29)))*(~(n57)))*(n489))))) ;
assign n2892 = ((n533)*(~((n193)*(n2884))))*(n4075) ;
assign n2897 = ((((n533)*(~((n193)*(n2884))))*(~(n1513)))*(n2317))*(n2892) ;
assign n4084 = (~(((((~(n6))*(~(n2207)))*(n2251))*(n2320))*(~(n2897))))*(~(n1504)) ;
assign n2911 = ((~((~(((~(n54))*(~(n55)))*(~(n56))))*(~(((~(n54))*(n55))*(~(n56))))))*(n79))*(n1311) ;
assign n2915 = ((((~((~(n487))*(~(n489))))*(~(n499)))*(~(n1311)))*(n1586))*(~(n2424)) ;
assign n2917 = (n151)*(~((n5)*(n2306))) ;
assign n4102 = ((((~((~(n81))*(n591)))*(~(n178)))*(n200))*(~(n1304)))*(~(n1311)) ;
assign n2975 = (~((~(n204))*(n205)))*(~((n204)*(~(n205)))) ;
assign n4109 = (~((((~(n54))*(~(n55)))*(~(n56)))*((n204)*(~(n205)))))*(~((n485)*((n204)*(~(n205))))) ;
assign n3056 = (n5)*(n2277) ;
assign n4116 = (~((((~(n204))*(n205))*(n206))*(~(n216))))*(~((n5)*(n2307))) ;
assign n3102 = (n46)*(n47) ;
assign n3103 = (n48)*((n46)*(n47)) ;
assign V321(2) = (~(((~((~((~(n578))*((~(n577))*(~(n578)))))*(~((n578)*((n578)*(~(n587)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n148))*(~(n661))));
assign V356 = (((((~(n1001))*(~(n1086)))*(~(n1114)))*(~(n1131)))*(~(n1148)))*(n3314);
assign V357 = (((((~(n1190))*(~(n1212)))*(~(n1235)))*(~(n1252)))*(~(n1269)))*(n3372);
assign V373 = (n7)*(n8);
assign V375(0) = ~(((((~((n53)*(n71)))*(~((n32)*(n53))))*(~((n53)*(n149))))*(n3380))*(n3381));
assign V377 = (n10)*(~((~(n9))*(~((((n10)*(~(n59)))*(n60))*(n65)))));
assign V393(0) = ~(((~((((~(n13))*(n38))*(n1309))*(n1313)))*(~(((~(n13))*(n1313))*(n1414))))*(~(n1406)));
assign V398(0) = ~(((((~((n1304)*(n1313)))*(~(n21)))*(~(n1406)))*(n3465))*(n3466));
assign V410(0) = ~(((~((~((n5)*(~(n1431))))*(n3474)))*((~((~(n204))*(n205)))*(~((n204)*(n205)))))*(~(n1311)));
assign V423(0) = ~(((((~((n15)*(n628)))*(~(n1313)))*(~(n1435)))*(n3450))*(n3451));
assign V432 = ((((~((n40)*(n1313)))*(~((n1304)*(n1313))))*(~(n1454)))*(n3509))*(n3510);
assign V435(0) = ~((~(n1601))*(~(n1616)));
assign V500(0) = ~((~(n24))*(n151));
assign V508(0) = ~((~(n1626))*(n3535));
assign V511(0) = ~((~(n25))*(~((~(n21))*(n26))));
assign V512 = (((~((n251)*(~(n252))))*(~((~(n251))*(n252))))*(~((n249)*(~(n250)))))*(~((~(n249))*(n250)));
assign V527 = ((((~((n3539)*(n3540)))*(~(n21)))*(~(n22)))*(~(n1311)))*(~(n1586));
assign V537 = ((~(n17))*(n485))*(~(n883));
assign V538 = ((~(n17))*(n485))*(~(n823));
assign V539 = ((~(n17))*(n485))*(~(n907));
assign V540 = ((~(n17))*(n485))*(~(n713));
assign V541 = ((~(n17))*(n485))*(~(n1679));
assign V542 = ((~(n17))*(n485))*(~(n1702));
assign V543 = ((~(n17))*(n485))*(~(n1725));
assign V544 = ((~(n17))*(n485))*(~(n1751));
assign V545 = ((~(n17))*(n485))*(~(n1777));
assign V546 = ((~(n17))*(n485))*(~(n1803));
assign V547 = ((~(n17))*(n485))*(~(n1830));
assign V548 = ((~(n17))*(n485))*(~(n1854));
assign V572(9) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(~(n1401)))*(n1865)))*(~((((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(~(n120)))*(~(n1865)))));
assign V572(8) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(~(n1363)))*(n1865)))*(~((~(n1865))*(n3631))));
assign V572(7) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(~(n1382)))*(n1865)))*(~((~(n1865))*(n3638))));
assign V572(6) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n1920))))*(~(((~((~(n501))*(n538)))*(~(n1865)))*(n3650))));
assign V572(5) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n1954))))*(~(((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(n3666))));
assign V572(4) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n1989))))*(~((((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(~(n1865)))*(~(n1998)))));
assign V572(3) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n2043))))*(n3701));
assign V572(2) = ~((~(((((~((~(n501))*(n537)))*(~(n501)))*(n538))*(n1865))*(~(n2090))))*(n3725));
assign V572(1) = ~((~((~(n1865))*(n3733)))*(n3749));
assign V572(0) = ~((~(((~((~(n501))*(n537)))*(~((~(n501))*(n538))))*(n3753)))*(n3758));
assign V585(0) = ~V34(0);
assign V587 = (~(n34))*(~((~((~(n70))*(~(n77))))*(~((~(n549))*((~(n537))*(~(n538)))))));
assign V591(0) = ~((~(((~((~((~(n70))*(~(n77))))*(~((~(n549))*(n566)))))*(~(n34)))*(n35)))*(~(((~((~((~(n70))*(~(n77))))*(~((~(n549))*(n566)))))*(n34))*(~(n35)))));
assign V597(0) = ~((~(((~((~((~(n70))*(~(n77))))*(~(n567))))*(~((n34)*(n35))))*(n36)))*(~(((~((~((~(n70))*(~(n77))))*(~(n567))))*((n34)*(n35)))*(~(n36)))));
assign V603(0) = ~((~(((~((n36)*((n34)*(n35))))*(~((~(n501))*(~(n567)))))*(n37)))*(~((((n36)*((n34)*(n35)))*(~((~(n501))*(~(n567)))))*(~(n37)))));
assign V609(0) = ~((~(((~((n37)*((n36)*(n1307))))*(~((~(n501))*(~(n567)))))*(n38)))*(~((((n37)*((n36)*(n1307)))*(~((~(n501))*(~(n567)))))*(~(n38)))));
assign V620 = (~((((~((~(n631))*(~(n1620))))*(n16))*(~(n22)))*(~(n1311))))*(n3775);
assign V621 = (n39)*((~((~(n26))*(n253)))*(~((n26)*(~(n253)))));
assign V630 = ((~(((~((n5)*(n598)))*(~(n41)))*(n3523)))*(~((n15)*(n598))))*(~(n40));
assign V634(0) = (~((n43)*((~(n24))*(~(((~(n24))*(n43))*(~(n44)))))))*(~(((~(((~(n24))*(n43))*(~(n44))))*(n24))*(n42)));
assign V640(0) = ~((~(n24))*(~(((~(n24))*(n43))*(~(n44)))));
assign V657 = ~V257(7);
assign V707 = (~(n57))*((~(n17))*(((~(n54))*(~(n55)))*(~(n56))));
assign V763 = ((((~((~(n485))*(n3159)))*(n69))*(~(n183)))*(~(n184)))*(~(n509));
assign V775 = ((((n20)*(n151))*(n513))*(~(n533)))*(n2254);
assign V778 = (n53)*(n71);
assign V779 = (n72)*((n7)*(~(n8)));
assign V780 = (n53)*(n72);
assign V781 = ((~((~(n70))*(~((~(n17))*((n5)*(~(n500)))))))*(n72))*(n73);
assign V782 = (n32)*((n7)*(~(n8)));
assign V783 = (n71)*(n74);
assign V784 = (n32)*(n74);
assign V787 = (n32)*(n53);
assign V789 = ((~(((~(n8))*(n44))*(n182)))*(n53))*(n75);
assign V798(0) = ~(((((~(n40))*(n151))*(~(n2298)))*(n2336))*(n3837));
assign V801 = (n500)*(((((n20)*(~(n61)))*(~(n62)))*(~(n63)))*(n76));
assign V802(0) = ~((~(n70))*(~(n77)));
assign V821(0) = ~((~((~(n80))*(~((~((~(n70))*(~(n77))))*((n57)*(n544))))))*(~((n29)*((~((~(n70))*(~(n77))))*((n57)*(n544))))));
assign V826(0) = ~(((~(((~((~(n501))*((n57)*(n544))))*(n80))*(n81)))*(~((~(n81))*((~(n80))*(~((~(n501))*((n57)*(n544))))))))*(~((n30)*((~(n501))*((n57)*(n544))))));
assign V966 = ((~((~((~((~(n70))*(~(n77))))*(~(n2298))))*(n3851)))*(n151))*(n2254);
assign V986 = ((~(((~((n15)*(~(n534))))*(~(n2366)))*(~(n2369))))*(n151))*(n2254);
assign V1213(11) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1840)))))*(~((n578)*((n578)*(~(n1846)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n136))*(~(n661)))));
assign V1213(10) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1816)))))*(~((n578)*((n578)*(~(n1822)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n137))*(~(n661)))));
assign V1213(9) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1790)))))*(~(n1797))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n138))*(~(n661)))));
assign V1213(8) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1764)))))*(~(n1771))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n131))*(~(n661)))));
assign V1213(7) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1738)))))*(~(n1745))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n132))*(~(n661)))));
assign V1213(6) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1715)))))*(~((n578)*((n578)*(n583))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n133))*(~(n661)))));
assign V1213(5) = ~((~(((~((~((~(n578))*((~(n578))*(~(n1692)))))*(~((n578)*((n578)*(~(n583)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n134))*(~(n661)))));
assign V1213(4) = ~((~((((~((n513)*(n534)))*(~((~(n593))*(~(n661)))))*(n661))*(~(n1672))))*(~((((~(n593))*(~(n661)))*(n135))*(~(n661)))));
assign V1213(3) = ~((~((((~((~(n593))*(~(n661))))*(n661))*(~(n703)))*(n3222)))*(~((((~(n593))*(~(n661)))*(n4))*(~(n661)))));
assign V1213(2) = ~((~((((~((~(n593))*(~(n661))))*(n661))*(~(n898)))*(n3252)))*(~((((~(n593))*(~(n661)))*(n3))*(~(n661)))));
assign V1213(1) = ~((~((((~((~(n593))*(~(n661))))*(n661))*(~(n814)))*(n3232)))*(~((((~(n593))*(~(n661)))*(n2))*(~(n661)))));
assign V1213(0) = ~((~((((~((~(n593))*(~(n661))))*(n661))*(~(n874)))*(n3242)))*(~((((~(n593))*(~(n661)))*(n1))*(~(n661)))));
assign V1243(9) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1396))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n139))*(~(n661)))));
assign V1243(8) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1358))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n140))*(~(n661)))));
assign V1243(7) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1377))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n141))*(~(n661)))));
assign V1243(6) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1915))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n142))*(~(n661)))));
assign V1243(5) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1949))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n143))*(~(n661)))));
assign V1243(4) = ~((~(((~((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661))))*(n661))*(~(n1984))))*(~((((~((n164)*(~((~(n538))*(~(n591))))))*(~(n661)))*(n144))*(~(n661)))));
assign V1243(3) = ~((~(((~((~(n593))*(~(n661))))*(n661))*(~(n2038))))*(~((((~(n593))*(~(n661)))*(n145))*(~(n661)))));
assign V1243(2) = ~((~(((~((~(n593))*(~(n661))))*(n661))*(~(n2085))))*(~((((~(n593))*(~(n661)))*(n146))*(~(n661)))));
assign V1243(1) = ~((~(((~((~(n593))*(~(n661))))*(n661))*(~(n2133))))*(~((((~(n593))*(~(n661)))*(n147))*(~(n661)))));
assign V1243(0) = ~((~(((~((~((~(n578))*((~(n577))*(~(n578)))))*(~((n578)*((n578)*(~(n587)))))))*(~((~(n593))*(~(n661)))))*(n661)))*(~((((~(n593))*(~(n661)))*(n148))*(~(n661)))));
assign V1256 = (n149)*((n7)*(~(n8)));
assign V1257 = ((((~(n9))*(~(n17)))*(n73))*(n149))*(n3868);
assign V1258 = (n53)*(n149);
assign V1259 = (n53)*(n150);
assign V1260 = (n74)*(n150);
assign V1261 = (~(n15))*((n74)*(n150));
assign V1262 = (n75)*((n7)*(~(n8)));
assign V1263 = (n53)*(n75);
assign V1264 = (n73)*(n75);
assign V1265 = (n70)*((n73)*(n75));
assign V1266 = (n74)*(n75);
assign V1267 = (n74)*(n149);
assign V1274(0) = ~((~((((n627)*(n630))*((n151)*(n2254)))*(n15)))*(~(n2413)));
assign V1281(0) = ~((~((((n151)*(~((n5)*(n2308))))*(n152))*(n2430)))*(~((~(n2430))*((~(n2430))*(~(n2439))))));
assign V1297(4) = ~((~((((n151)*(~((n5)*(n2308))))*(n153))*(~(n2429))))*(~((n2429)*((n64)*(n2429)))));
assign V1297(3) = ~((~((((n151)*(~((n5)*(n2308))))*(n154))*(~(n2429))))*(~((n2429)*((n63)*(n2429)))));
assign V1297(2) = ~((~((((n151)*(~((n5)*(n2308))))*(n155))*(~(n2429))))*(~((n2429)*((n62)*(n2429)))));
assign V1297(1) = ~((~((((n151)*(~((n5)*(n2308))))*(n156))*(~(n2429))))*(~((n2429)*((n61)*(n2429)))));
assign V1297(0) = ~((~((((n151)*(~((n5)*(n2308))))*(n157))*(~(n2429))))*(~((n2429)*((n76)*(n2429)))));
assign V1365 = ((((~(n1514))*(n2397))*(n534))*(n647))*(n3911);
assign V1375 = ~V268(5);
assign V1378 = ((n32)*((n7)*(~(n8))))*((~(n501))*(~((~(n537))*(~(n538)))));
assign V1380 = (n2266)*(~(((~((~(n566))*(n3922)))*(~((~(n1858))*(n3927))))*(~(n1864))));
assign V1382 = ((~((~(n591))*(~((~(n501))*(~(n1580))))))*((n7)*(~(n8))))*(n32);
assign V1384 = (((((n5)*(n32))*(~(n1311)))*(n1576))*(~(n1584)))*(n2259);
assign V1386 = (((~((~(n193))*(n533)))*(~(n2508)))*((n7)*(~(n8))))*(n32);
assign V1387 = (n53)*(n163);
assign V1392(0) = ~((~((n2397)*(n3942)))*(~((((n78)*(~(n628)))*(~(n1513)))*(n2397))));
assign V1423 = (n31)*(n53);
assign V1426 = (n31)*((n7)*(~(n8)));
assign V1428 = (n31)*(n74);
assign V1429 = (n31)*(n73);
assign V1431 = (~((~(n8))*(n167)))*((n31)*(n53));
assign V1432 = (((((~(n40))*(~(n1457)))*(~(n2207)))*(n2251))*(n19))*(n151);
assign V1439(0) = ~((~((~(n28))*((n30)*(n492))))*(~(((n151)*(n168))*(~(n538)))));
assign V1440(0) = ~((n151)*(~((n169)*(~((n168)*((~(n17))*(n485)))))));
assign V1451(0) = ~((~((((~(n2509))*(~(n2535)))*(n85))*(n151)))*(~(((~((~(n2509))*(~(n2535))))*(~(n85)))*(n151))));
assign V1459(0) = ~((~((((~((~(n85))*(n2509)))*(~((n85)*(n2535))))*(n151))*(n170)))*(~(((~((~((~(n85))*(n2509)))*(~((n85)*(n2535)))))*(n151))*(~(n170)))));
assign V1467(0) = ~((~((((~((~(n170))*((~(n85))*(n2509))))*(~((n170)*((n85)*(n2535)))))*(n151))*(n171)))*(~(((~((~((~(n170))*((~(n85))*(n2509))))*(~((n170)*((n85)*(n2535))))))*(n151))*(~(n171)))));
assign V1470 = (((~((n28)*((~(n30))*(n596))))*(n151))*(n172))*(n2254);
assign V1480(0) = ~(((~(((~((~(n70))*(~(n77))))*(~((~((~(n204))*(n205)))*(~((n204)*(n205))))))*(n544)))*(~((~(n544))*(~((~((~(n204))*(n205)))*(~((n204)*(n205))))))))*(~(n1584)));
assign V1481(0) = ~V214(0);
assign V1492(0) = ~((~((~(n22))*(n175)))*(~(((n18)*(n151))*(n3956))));
assign V1495(0) = ~V175(0);
assign V1512(3) = ~((~((n2251)*(~(n2591))))*(~((n2591)*(~((((~(n1235))*(~(n1252)))*(~(n1269)))*(n3979))))));
assign V1512(2) = ~((~((~(n2591))*(~(n2603))))*(~((n2591)*(~((((~(n1148))*(~(n1207)))*(~(n1235)))*(n3988))))));
assign V1512(1) = ~((~((~(n2591))*(~((n2251)*(n2261)))))*(~((n2591)*(~(((~(n1190))*(~(n1252)))*(n3997))))));
assign V1536(0) = ~((((~((n544)*(n1586)))*(~(((n5)*(n27))*(n544))))*(n2251))*(~(n2585)));
assign V1537 = (((((~(n40))*(~(n1457)))*(~(n2207)))*(n2251))*(n151))*(n173);
assign V1539 = ((~((~(n174))*(~(n180))))*(n151))*(n2254);
assign V1552(1) = ~((~((((~((~(n501))*(~(n1580))))*(~(n110)))*(n501))*(n591)))*(~((((~(n501))*(~(n1580)))*(~((n501)*(n591))))*(~(n1401)))));
assign V1552(0) = ~((~((((~((~(n501))*(~(n1580))))*(~((~((n110)*(~(n111))))*(~((~(n110))*(n111))))))*(n501))*(n591)))*(~((((~(n501))*(~(n1580)))*(~((n501)*(n591))))*(~(n1363)))));
assign V1613(0) = (~((~((~((~(n2657))*((~((~(n2671))*(n2690)))*(~((n2671)*(~(n2690)))))))*(~((n2657)*(~((~((~(n2671))*(n2690)))*(~((n2671)*(~(n2690))))))))))*(n2781)))*(~(((~((~(n2657))*((~((~(n2671))*(n2690)))*(~((n2671)*(~(n2690)))))))*(~((n2657)*(~((~((~(n2671))*(n2690)))*(~((n2671)*(~(n2690)))))))))*(~(n2781))));
assign V1613(1) = (~((~((~((~(n2797))*((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))*(~((n2797)*(~((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811))))))))))*((~((~((~((~(n2824))*(n2831)))*(~((n2824)*(~(n2831))))))*(n2851)))*(~(((~((~(n2824))*(n2831)))*(~((n2824)*(~(n2831)))))*(~(n2851)))))))*(~(((~((~(n2797))*((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))*(~((n2797)*(~((~((~(n2804))*(n2811)))*(~((n2804)*(~(n2811)))))))))*(~((~((~((~((~(n2824))*(n2831)))*(~((n2824)*(~(n2831))))))*(n2851)))*(~(((~((~(n2824))*(n2831)))*(~((n2824)*(~(n2831)))))*(~(n2851))))))));
assign V1620(0) = ~((((~((n17)*(n1311)))*(~((~(n40))*(n183))))*(~((n17)*(~(n2251)))))*(~(n509)));
assign V1629(0) = ~(((~(((~(n187))*(~(n1513)))*(~(n1620))))*((~((~(n26))*(n253)))*(~((n26)*(~(n253))))))*(~(n2867)));
assign V1645(0) = ~(((~((n27)*((~((~(n70))*(~(n77))))*(n544))))*(~(n1523)))*(~(n2424)));
assign V1652(0) = ~((((((~(n193))*(n533))*(~(n14)))*(~(n79)))*(n189))*(n4069));
assign V1669 = ((~(((~(n6))*(~(n2328)))*(n2892)))*(~((n501)*((~(n6))*(n1457)))))*(n4084);
assign V1671(0) = ~V205(0);
assign V1679(0) = ~((n533)*(~(n2884)));
assign V1693(0) = ~((~((((~(n2911))*(~(n2915)))*(n194))*(n2917)))*(~((~((~(n2911))*(~(n2915))))*((~(n2439))*(~((~(n2911))*(~(n2915))))))));
assign V1709(4) = ~((~((((n151)*(~((n5)*(n2306))))*(n195))*(~(n2911))))*(~((n2911)*((n64)*(n2911)))));
assign V1709(3) = ~((~((((n151)*(~((n5)*(n2306))))*(n196))*(~(n2911))))*(~((n2911)*((n63)*(n2911)))));
assign V1709(2) = ~((~((((n151)*(~((n5)*(n2306))))*(n197))*(~(n2911))))*(~((n2911)*((n62)*(n2911)))));
assign V1709(1) = ~((~((((n151)*(~((n5)*(n2306))))*(n198))*(~(n2911))))*(~((n2911)*((n61)*(n2911)))));
assign V1709(0) = ~((~((((n151)*(~((n5)*(n2306))))*(n199))*(~(n2911))))*(~((n2911)*((n76)*(n2911)))));
assign V1717(0) = ~((~((n2254)*(n4102)))*(~((~(n501))*(~((~(n591))*(~((~(n540))*(~(n567)))))))));
assign V1719 = ((~(((n59)*(~(n60)))*(n65)))*(~(n178)))*(n200);
assign V1726(0) = ~((~(((n151)*(n201))*(n566)))*(~(((~(n567))*(n1858))*(n2591))));
assign V1736 = ((((~(n6))*((~(n64))*(n1311)))*(~(n79)))*(n501))*(n1604);
assign V1741(0) = ~(((((~((~(n1311))*(n2219)))*(~((n79)*(n1311))))*(~((~(n1311))*(n2225))))*(~((~(n1311))*(n2228))))*(~(n2216)));
assign V1745(0) = ~((((n6)*(n203))*(~(n485)))*(~(n499)));
assign V1757(0) = ~((~((~(n204))*(n205)))*(~((n204)*(n205))));
assign V1758(0) = ~((~((~(n204))*(n205)))*(~((n204)*(~(n205)))));
assign V1759(0) = ~((~(((~((n5)*(n2278)))*(n151))*(n206)))*(n4109));
assign V1760(0) = ~V101(0);
assign V1771(1) = ~((~((n598)*((~(n67))*(n598))))*(~((~(n598))*((~(n244))*(~(n598))))));
assign V1771(0) = ~((~((n598)*((~(n66))*(n598))))*(~((~(n598))*((~(n245))*(~(n598))))));
assign V1781(1) = ~((~((~(n598))*((~(n598))*(n1854))))*(~((n598)*((~(n248))*(n598)))));
assign V1781(0) = ~((~((~(n598))*((~(n598))*(n1830))))*(~((n598)*((~(n247))*(n598)))));
assign V1829(9) = ~((~((n23)*((n23)*(n1401))))*(~((~(n23))*((~(n23))*(n667)))));
assign V1829(8) = ~((~((n23)*((n23)*(n1363))))*(~((~(n23))*((~(n23))*(n1854)))));
assign V1829(7) = ~((~((n23)*((n23)*(n1382))))*(~((~(n23))*((~(n23))*(n1830)))));
assign V1829(6) = ~((~((n23)*((n23)*(n1920))))*(~((~(n23))*((~(n23))*(n1803)))));
assign V1829(5) = ~((~((n23)*((n23)*(n1954))))*(~((~(n23))*((~(n23))*(n1777)))));
assign V1829(4) = ~((~((n23)*((n23)*(n1989))))*(~((~(n23))*((~(n23))*(n1751)))));
assign V1829(3) = ~((~((n23)*((n23)*(n2043))))*(~((~(n23))*((~(n23))*(n1725)))));
assign V1829(2) = ~((~((n23)*((n23)*(n2090))))*(~((~(n23))*((~(n23))*(n1702)))));
assign V1829(1) = ~((~((n23)*((n23)*(n2138))))*(~((~(n23))*((~(n23))*(n1679)))));
assign V1829(0) = ~((~((~(n23))*((~(n23))*(n667))))*(~((n23)*((n23)*(n907)))));
assign V1832 = (n151)*(~((~(n2535))*(~((n192)*(~(((n193)*(~(n2508)))*(~(n2884))))))));
assign V1833(0) = ~V261(0);
assign V1863(0) = ~V301(0);
assign V1864(0) = ~V302(0);
assign V1896(0) = ~(((~((n212)*(~((n5)*(n2277)))))*(~((n204)*(n205))))*(~(n1584)));
assign V1897(0) = ~((~(((~(n17))*(n485))*(n1584)))*(~((n213)*(~((n5)*(n2277))))));
assign V1898(0) = ~((~((n485)*(((n18)*(n172))*(n178))))*(~((n214)*(~(n3056)))));
assign V1899(0) = ~((~((n487)*(((n18)*(n172))*(n178))))*(~((n215)*(~(n3056)))));
assign V1900(0) = ~((~((~(n204))*(n205)))*(~((n216)*(~((n5)*(n2277))))));
assign V1901(0) = ~((~((n204)*(~(n205))))*(~((n217)*(~((n5)*(n2278))))));
assign V1921(5) = ~((~(((((n218)*(~(n2277)))*(n2301))*(~(n2306)))*(~(n2308))))*(n4010));
assign V1921(4) = ~((n4017)*(n4018));
assign V1921(3) = ~((n4023)*(n4024));
assign V1921(2) = ~((n4029)*(n4030));
assign V1921(1) = ~((n4035)*(n4036));
assign V1921(0) = ~((n4041)*(n4042));
assign V1953(1) = (((n230)*(~(n2278)))*(n2301))*(~(n2307));
assign V1953(7) = ~((~((((n224)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n232)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(6) = ~((~((((n225)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n233)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(5) = ~((~((((n226)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n234)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(4) = ~((~((((n227)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n235)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(3) = ~((~((((n228)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n236)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(2) = ~((~((((n229)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n237)*(~(n2278)))*(~(n2301)))*(n2307))));
assign V1953(0) = ~((~((((n231)*(~(n2278)))*(n2301))*(~(n2307))))*(~((((n217)*(n2278))*(~(n2301)))*(~(n2307)))));
assign V1960(1) = ~((~(((n238)*(n1628))*(n2307)))*(~(((n240)*(~(n1628)))*(~(n2307)))));
assign V1960(0) = ~((~(((n239)*(n1628))*(n2307)))*(~(((n241)*(~(n1628)))*(~(n2307)))));
assign V1968(0) = ~((~(((n151)*(n243))*(n4116)))*(~(((~((~(n242))*(n2975)))*(~(n243)))*(n487))));
assign V1992(1) = ~((~((((~((~(n1860))*(~((~(n501))*(~(n566))))))*(~((~(n501))*(~(n566)))))*(~(n244)))*(n1860)))*(~((((~((n1860)*(~((~(n501))*(~(n566))))))*(~((~(n501))*(~(n566)))))*(n244))*(~(n1860)))));
assign V1992(0) = ~((~((((~((~(n1860))*(~((~(n501))*(~(n566))))))*(~((~(n501))*(~(n566)))))*(~((~((n244)*(~(n245))))*(~((~(n244))*(n245))))))*(n1860)))*(~((((~((n1860)*(~((~(n501))*(~(n566))))))*(~((~(n501))*(~(n566)))))*(n245))*(~(n1860)))));
assign V650 = ~((~((n130)*(~(((((n49)*(n50))*(n51))*(n52))*(n3103)))))*(~((~(n130))*(((((n49)*(n50))*(n51))*(n52))*(n3103)))));
assign V651 = ~((~((n49)*(~(((((n48)*(n3102))*(n50))*(n51))*(n52)))))*(~((~(n49))*(((((n48)*(n3102))*(n50))*(n51))*(n52)))));
assign V652 = ~((~((n50)*(~((((n48)*((n46)*(n47)))*(n51))*(n52)))))*(~((~(n50))*((((n48)*((n46)*(n47)))*(n51))*(n52)))));
assign V653 = ~((~((n48)*(~((((n46)*(n47))*(n51))*(n52)))))*(~((~(n48))*((((n46)*(n47))*(n51))*(n52)))));
assign V654 = ~((~((n51)*(~((n52)*((n46)*(n47))))))*(~((~(n51))*((n52)*((n46)*(n47))))));
assign V655 = ~((~((n47)*(~((n46)*(n52)))))*(~((~(n47))*((n46)*(n52)))));
assign V656 = ~((~((~(n46))*(n52)))*(~((n46)*(~(n52)))));
assign V1370 = ~((~((n207)*(~(((((n158)*(n159))*(n160))*(n161))*(n162)))))*(~((~(n207))*(((((n158)*(n159))*(n160))*(n161))*(n162)))));
assign V1371 = ~((~((n160)*(~((((n158)*(n159))*(n161))*(n162)))))*(~((~(n160))*((((n158)*(n159))*(n161))*(n162)))));
assign V1372 = ~((~((n161)*(~((n162)*((n158)*(n159))))))*(~((~(n161))*((n162)*((n158)*(n159))))));
assign V1373 = ~((~((n159)*(~((n158)*(n162)))))*(~((~(n159))*((n158)*(n162)))));
assign V1374 = ~((~((~(n158))*(n162)))*(~((n158)*(~(n162)))));
endmodule

